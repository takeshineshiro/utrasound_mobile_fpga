// megafunction wizard: %LPM_ABS%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_abs 

// ============================================================
// File Name: ABS.v
// Megafunction Name(s):
// 			lpm_abs
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.0 Build 132 02/25/2009 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module ABS (
	data,
	result);

	input	[29:0]  data;
	output	[29:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: OptionalOverflowOutput NUMERIC "0"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: nBit NUMERIC "30"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_ABS"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "30"
// Retrieval info: USED_PORT: data 0 0 30 0 INPUT NODEFVAL data[29..0]
// Retrieval info: USED_PORT: result 0 0 30 0 OUTPUT NODEFVAL result[29..0]
// Retrieval info: CONNECT: @data 0 0 30 0 data 0 0 30 0
// Retrieval info: CONNECT: result 0 0 30 0 @result 0 0 30 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL ABS.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ABS.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ABS.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ABS.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ABS_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ABS_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
