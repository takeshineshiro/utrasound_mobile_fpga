��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω����	8��7���I�N<��;���Z��4d��{�
��|��Ȋ)zo1���á�K���b��j.~���m��+?��bV��ݙ���M7\F���r��C>C�݂�N$��/���	�0���'v6�o�*�HA6�Ѡ��s-�v��x�۔7�D��:�b�#�Bn�K�͎��uP!ߌ��˼�{�&��t�7H��'jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��V�)��[�P��;�� 9�/�<"����_quf�tg����_��9(?��lds£����&��^z[��K�j��c�*z�w4G� ���������	x]̍��;��7�I��"8YdK�o����Oh5��&}Xa��gR�ca������pN�Wu��w)�S��X3����~篟|��ᕧSt ��[֊��Jџ�_�v%䆘[m�~R���\D�	m�!=�y����h�}�)���32�)���K��OC���N^o?�M��;]���i͹�9 ���t��%���&Oǀ�Һ�3{����V���	x]�<���eQ���X��\���|�@c���Կ�:�%n��e�ι̕��R)U�~�O���`Y�5���=�zX4P?�o��ľ��UW��͌Tfu��w)�S �J���vy7��Mv�9�h�s����b�z�Y8�:r&@�	��Ϸ)�����V\~{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�T�`�7?�\��4�/�I����D;�~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/�R����+��T��D[I'�p\���nEA���KW\�#Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hG[��{�ĘX�������_�~/�F߼
�dr���3/7D�d�/+M���"��ei,l����Fv!.�僢�#��i����S(�Z���kv
�u��7+�����I�>g���#�W�w��fD�5����`K�P�C�s�&R�߷�C�Q���clׇ��I�����o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��g�,P�ny�ӓ���&D�H��V�6IWJE�r���秹��ч��~3�V0U�	�I]���T���u�If:i�!��B���y�4r7h��Ϭ�c�8(;��w��!�+�7����ݸb��3���ne��'�{�a����'3��n��W�߼
�dջ{5NHdY��~<��Q�5}�m�0��o��7�ܥ��2�nhτ���ˈ�s������2]N�X�cdA!���o�I�?g�fY�~�a���+�Uz�QL���}�'����"�|�E+��T��D[I'�p\���nEA�_42K2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��ݞƼ�FmEOН9_l8K,H"��sD�sK~,�t,X�0��y>@���D��!r �z�듻�D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��}�`wKݷ/���W�8yQ�5}�m�0��o��7�ܥ��2�nhτ���ˈ�s������XP��~�26��\��Y���eʆ�In��t��+x�r�u�#��nt��c�s5jݭ�F����μ<�e<�^��XzHL� ��C�7ª6��O��/$Z��Qu���%$��>_��̃x0�?��t�7h���;�jmT�#~�ty�#�"��dѓ�u��r��Ƹv��*QxR��9�H�@�}S�L�#�x�첎Ϡp�bO(�����/�x�첎���K�N]�H&� �!�`�(i3�q{�).+95���g�֕�0N�s2fĉ>99��A0ok�?�JY�)�Y`��jD4��S��c��څH�8��)<��U��tT��kU�t���o�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����47��"(;�8���%7)��۟�08ݭ�Q<���2�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX��W<���ubr�N���,�ƺ =�Uvc�8(;��w��!�+�7����ݸb��3���ne��'�{�a����'3:{%:k�a�2N��n�âW[��8u�n�B��t�t>
xL�Q�S�ֱ�q�����)�@t(��֚��\�v�M��%�p@��=H��F�Z�B? M�7FG��P�v�"�L���n3�ڌybN}�m��{�!����� V�"����Q�)�@�ֱ�q������m�q�)Ў6dG��O����14�7'U�1sly�d2N#�8&���I���A��y�u���1ИdN�<@Iv�O�ȕi�g}|�H�q�M'�y���~+�ݗ7�%M���y�(0��7��ZX#(� �301�f�[��(����#�a�Ą�[�J�iP]m��m�H�RtV�^C��r��Si	F�������,�˞��X��/��e]t�ˇ�ۅ"0�ď�B�'��a�q�M'�y���~+�ݗ�"�чE4����k[J@&�4�T�TN���K�Ǔ�\u���1ИdN�<@Iv�O�ȕi��:5A��p��jVѭ@�K�Ǔ�\��ub-���8�-5
�h|L8�~���@�VҒm͢����z��Q�ye�M�8pƣ��  6 y2��R���Ě����E�i�m}640�RS���$
�)��A�?�j�#���y��5Sà�+�\b��5M2Wŀ;s���}(ʥ�nr]�b�N���UsMDZK� j��������n7,�ڻC�i��9���1�L�]�b�֘m��+?��bV����
~�d�!N�'�y�G