��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9|[�,HJ
Κ�P/�u�x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`��;�É_g�?�H�.J"����U���T���딣0&_���X0���2|	p��rw@	@us��n��/�FI���O8�yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|�o�r� �K�����)�݉|�7\F���r��RL�a)ѻtUWR����H7��7�ޑ����<��&g�7C��H��C=�)3�C����")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|?_W�\I��^�َ2V�N�u�k1i�f1?�نN��_�Q�L���E�aC�h�>�N{a�9O��Yk"1/>���M[�a7Y��0�-�R$��Ct�z&��ÃlO ܅dh�' L� U��֜��3jݭ�F���L�D��6S�]V�H7'�R�^Ƒ���a�\����9�	��%т��!o.sG[�� �`�>:8�A�/����<.+6J!�t���\�W��F�eD4];ˍH�7��_��T��!e����\G�YIpsl�ć���vh�ҋX������S8�J�]=��R�^Ƒ����"X��[��Q[R�7�%=��L�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y����q��G8�����b,�e.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7&�e��A�����
L'���Xw�j�7��ct�:��RE��W��_�ړ8���/��4��}�<�e�y���J�@IE�U����S8�/ #O�)R�^Ƒ����"X��[�d�a�4$��9+�����o��C!T*�q���U����?�N�By3��<Z鎬�����X���*_��(֥�S�)37J*u>����CΫa������<��z��}���w�V�"-4��h�]8+��T����oGo�Z�K����ހ d�����L��]�>-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/>���M[�a7Y��0�-�R$��;g��4��s;�s��&<�w�п?G��q8h�G[�� 4&Ƒ:2�c<�^<�H�U�YQN`V��	��y��2����8��`+S6E���7-K����}�)��E�d�-���geW���w>��Y��$1&ODQ3�z�sis@�����]���ϸ��#|S������3[�u8�J�a3mPy��>/' k!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�����hWK{m35%7� ��yDg!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����hWK{m35%,�!�H<�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����h�? "a��Q�V!�(�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�����h�? "a��%}w�dN�!�`�(i3�X;p`�V�׍A�f�?ǉ�=�t� ��O���}���i!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�$�V��bst�N���!�`�(i3!�`�(i3�X;p`���z�����2� ��=�<���� z!�`�(i3!�`�(i3!�`�(i3�sg]�_�}F�r�f�t��5Z�����N���96!�`�(i3!�`�(i3!�`�(i3���I�=|�0��E|�,���6%�az\�m���Iϕ������z_۬=�!�`�(i3�&8�,�g����=�'�j���#�|M�d�>b�eIG��Q�q>x�-#F\eڲ!�`�(i3!�`�(i3��g��E��� ������$Y� 2��4�b��{�P}�!�`�(i3!�`�(i3�b[�u2�G�=����ڄ���������622���k˗S�d�!�`�(i3!�`�(i3@�C,��ǣ©��S:H��+܆} �S�
â!�`�(i3!�`�(i3-���d	c�b�ǣ©��S:H��+܆��K����!�`�(i3!�`�(i3-���d	c�b�ǣ©���_`Ogkl@`��m'��r�Nt[NzigzA=v)-��,ufOX�mCf�?ǉ�=�$Nx���t��y(�����������(����������)��-�L�߯d�8a,�X����>[H��_0Vձ!�`�(i3!�`�(i3�&8�,�I���Ut�es��O!�`�(i3�N�v�1��B�r��!�`�(i3!�`�(i3�$wq�����0��E|�,���6%�a����>[HÛON�?��!�`�(i3!�`�(i3�&8�,��w�Iſ�Κes��O!�`�(i3k�-i�9~�!�`�(i3!�`�(i3!�`�(i3�u~xgA���������6%�a����>[Hs�?����H�Ud���7!�`�(i3�&8�,�|�1�0j�~�Y���(���8���VZ��W�d�!�`�(i3!�`�(i3��5�q	�`
 ֢����e���W�\�h��&2��>/' k!�`�(i3P*N�2���9�����޲�e S]#�e����kn4@Q�/�!�`�(i3n&����_�a�/!O�f�?ǉ�=��9K��r|%oO���m�
��,!\4L$ֵ���A��)}�����*��hy�t�]�|����*[UxG!�`�(i3N>�X�5G���oy���ݚ�Н��@����MTl�������l6��6�5�p��`�T1)��/Z鎬�������(����z?|��f�?ǉ�=J�a3mPy�D`}Q'���Xw�j�7���z��0��ݚ�Н���O�q�̍YY~����V�my$�N�m��y���wӨj]h��0kI��h��d�)bU/�'5���ĭ�*�����X;p`�Z����c!�`�(i3�%]�N����%ў׫�t�$��o؍��R��w�R���y_Nr`e���4)���>݈��K+:��0	��