��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�յ�'�)���Ҷt������5O|�7x��������&�ǝ�+zA��]��~ا@H;�W ��W�5�k�s����F��W��`��q�©���?��P>����M7\F���r��C>C�݂�N$��/���	�0���'v6�o�*�HA6�Ѡ��s-�v��x�۔7�D��:�b�#�Bn�K�͎��uP!ߌ��˼�{�&���7�os!w����]��4�:j�l�,9����=-��Ǘ��p��W*[��HMiL���om�Q*���T�K�MV}xj\�iW�(� 0�D�A~����p��ؚ�fD�~����pn��-�4ڭ	���
��M!�nz��m��+ r���7�����|�]��;�I�Qg�@zh�S҆�|n����Շ_ Q -���W}�+��X��J�Й�m����u�����w`q�tc�ؑ��g�=Iĩ�m��d�7�Q����.P2:}��>�,�_'�hQr�k@Q��j��C�뫰v]uR����Pl����N�Er��xXc)O�%���ʅ�$n��RL�a)=�y�~ ���G�/9��i�:��^��I��X�7C��H���j�v�?�*�u��q[o��>�`u^9�렕4��S��$[��������\�4�sP	�b\qB��������"^Y怄�GW���և~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��ED�D ���
r:�����u��w)�S�5� �7��Mv�9*���f��^(��f�)y�8�:r&@��=��$얃�rb2 �Q[1I�����w'�\�Q�3M���e�t��yn�	� �x�m��n~�q({L�51��;����'��%Ճ�86���H�aF��6��I���j�r�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�E�s��bc�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�f{*n/�,傴����'SR����.�}|��ι%9M��j@�����nEAJ_�'��P9�tw:g+��T��٤�2[51g��f�PH2E���ƪϤ�Yk"1/��L�lW��+�va��2鍔�	g\A��AOge���ħƿ�9c�I�?g�f�$��P�`
5��*�z��Yk"1/���%	v3����M�}�O��ɝ�^�&d�A|?_W�\I���aC�h�>�N{a�9O��Yk"1/���]���l�uq9����ea�;y� ����t����M���������b9����4�6�t�����\{F˯�+)��n̈́�zL͊�q���Vǃ���߼��� .�����ݞ��D	��U����	�I	"k�+��v��z�N������i��b9����:ߐ�؍��R��j�.(Wx*��|��p��h�d �'���Xw�f�VHF��>BH<M�z�]�!����M[��Ǣ����K? T�ҋX����>��l%i�-"K��^��Hm��S�)37J*u�������ݹ�0����['����?���F��ʙ@E>*;�¬pX��g��U-�e�,���6+��\�!wn�Ŕ"�����/Z鎬����
C��8q��f�kN�ı��XK��(�W�~:n=�ct�:��RE��W��_�ړ8���/��4��}�<��/�^�Ӭ����
L'���Xw s4S�'�i��`�z��4�+|'Tԕ���ߋI7��-5|>����n�xY�J��ev�mS��0�-����#u��Yk"1/���]���lN��;
�'�����N<���d�k��Yu>�G Oag�qod�֓��+��T�����h�6ؖ� onc�9���$1m���/��&l�L��M�,���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7⏇���;�z*���Be�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)ƛ�>�֔�ټ*w2�56����n9�y2eŋU�sl�L��M�,���	N^�U{xN��i>r�<Uee�,��3�L��-+��B�G����n9�)��(��l�L��M�,���	N^�U{xN��i>r�<Uee�,��3�L��-+��B�G����n9�`�.E�y�ZWpH7���
I@1�ؠ&���Z02��`�z��4�+|'yG`ݜk��ʅ�-`[�=�5x�����c��D�of�7���A3�(N��㎏qló��@d��שt�v��I�`2ڻ�Ϊi3�|)sՀ�T:���V�Ra��l��!K��tf��
_�n�@/%{�;����f�kN�ı��XK��(ړ�8ݻ<�_���,D��{r81�ld�����WpH7���
I@1�ؠ&���Z02��`�z��4�+|'yG`ݜk�s��d�\��1+�v�[��P :��R'cf���³5����XK��(��s�Ӻ���?�d���&��ꢤ�Og0�oB��Z'N��;&�0z�cUL��,}w��kO��u����\�j��H���~���J��sa�"��q�Z鎬�������(���ܚ�2�E=hL�1p/-����#�p�t����M~V��	��y�����5�Dy�T^l;;��?:�e�{��x���#xW��z*K��t�v��I�`2ڻ�Ϊ;��|B���AW�*��G�J�����2wG!�'����ֈ|׸�F�5�O�%E#Pl�i�<�9��ݠ�.���?r$��Z鎬�������(���kO��u�}���	�f��/�Pqh.X �#_�惰�'�)�Բcf�b$j�p�t�v��I�`2ڻ�Ϊ���&3�{�H���~��w�R���y�\���_U�In��u��!�j��=)\�\��Eyz?]4��jyP����š��鶵��d���!i֭�h��O�׸��D������q��]�!��	Ǹ�y85�E���h�/	AT�D����$�P=Q�f}n�Z҇a,]v1�_ُ�}�Gv�['����?���F�- s
�VX7 �U6�.�g3Zdj�t���q��Sn(�JZ�Vk�;��|B�� �uR(ǜ`����ƫg�Tz�����;��|B����ҍ<��)#��!�&�kčw�⽒���M��������qb	��G��W+��W�}�t�sg6�o8:4�I���c�90�Ǘa��x[�����(����<m���"sS<�0�zG�������&G!�`�(i3��b`Һ�4	M+��I�}��nF���<�W�.�P�	��
�Q�}�߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3܌;���'����u��r��!�`�(i3��,� �݂��\���/Y��rx��"�@�����q ^C�Đ���%>�rGO�D mWN���%>�rGO�D mWNHN��R���IX0F�M��"����Y����,�ǰ�B`v���e?㙚7u6j�"Hs!���h5���kPc5��C�N�흰,_���9�+��O�r!�J��:�����lTN��IY��rx��"��9�ڮW;��|B��}��q4F�x�h�k�v�%�zq_҂T�q�w���t�v��I�`2ڻ�Ϊ_��s�֙R���Bk�d�C�JFɵ�&~����w�1&NXs;�¬pX��D�P�E6�k��q��־�W+��W��p����,D��������>���K�QZ���>�:5A��pCNZKE��e��#ɱ��\�!wn����t`x;��E�i�m}66j�"HsX�q&�^9Z���;��|B31F��~Gf��x��9�Mgw�� 
~�F�,���XF:��4�+|'\�����?�d���&��Xd��8�(J�yؕ�o!�'���4��Ǳ߁R�^Ƒ��D�P�E6�k��q��־�W+��W�2W���R0_.��45��LҺ_.E��p���V�$r�t�}iV��	��y�� �P�qN�/9ݦ�����,�ǰ� Ϳ�&�v��dY��0X2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��|�GJ Ւ�&�!x�� {k���o��W}d}��A�xm��ǯ+��3G�.��q�/@��۲�b�����A@�r$��E�V��Q"}Hi����k	���	5���n2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�3�n���SE`|Ň��O%��<�ν^Z�|Z��>B!�`�(i3 I���¬B���{�sc��ܯ�AZY��s��~!�`�(i3�% ���"�y&YA�%8�<Ŀ�]N�ұ|U
��4�5�ڜ���b��z�����p�_�/V��d��7�e��	t���3�q�Z�d�=��R"�磡�55�tץ���
��[H~��|vӥ{?�VU�簦!N�'�y�G