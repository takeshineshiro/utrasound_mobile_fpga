��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����i�'������\ᨅh��~�a.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I��7��?'�q�Z\�R�F*}Ø���K�Z�I�?g�f���\X�<����8��U�/?��qᾪ���>�*z�w4G�� ��d�n}K-J��K��z������3�z�ω���D���+��O����F72��{L�8br�.�/�d�������4�;���u�$|�>I��4�`���څk���ʬ~���t�켻�S���c,�8[0p����̀���1 T�V	�tL��	�<�A�}Q��"<�U���y�!u��&���.eԈ�{
��te�C��c�S+dk�%��G*)��L����R^�g�EP�O�.�A"V���2�uhǰv�%�]��I�uEd�=�>|(x������D�ԅ1Qr������i��Z��DN�n�������������8*��#�N�L~�4��,J�l�/���&�\ׇӭ��!�`�(i3!�`�(i3ɬc��WN������J��(<W]I� :��
&T������NUl��F�0?�R��e��/m
MN���q�p�8�s$%.F���=�Z&a_<t!�`�(i3!�`�(i3RaJ��te�.��vJw '��
�<s݌�����m�e6؟�r�Y�}94�h�z��/��PQ�A~}��/*0�(b��g��k���M���ʜ�Jo+{)�x�=�= s!�`�(i3!�`�(i3�J܏��٢���w���,ա�	r�?�#✲�@��1��A��'gKx/அ����`��o�)Wu�!�`�(i3!�`�(i3J�Y,�~)�{lN}Q�b�o�m�����m�e6��C�/�y9.Y'`f��������L�}��xİ k�ʞ�kĶ�r:w9���י�H[��e�ׇӭ��!�`�(i3!�`�(i3����n,��>]��e��2�qj�h�7pp����2u~-��)B�Kܓ!�`�(i3!�`�(i3��&'�y����s��.���Z�!Z��`�($+����������-N��]�1�l0�)�Myիnň��h����]ߺ�`@��h�h����M����CN�u!�`�(i3!�`�(i3��7���,�K�!5�����n,��'�\�n���t�u�?9Pjp��h���~��G����a�����(�I�?g�f���\X�<����8��U�/?��qᾪ���>�*z�w4G� ���������	x]��/$��x��~篟|�Q�M�u�cX8N_�=rџ�_�v%����E�)��|������\�4�sg�oXx��U������ՈĀO��w���9*<��*{�ۤ���*c���4�a6�N��?���\z-��EM���
+����rx�]�V��\#O���o�x��`�|>o}h5-*����>�xΕ���}�P�������pC-��h��☂/x+��s(a�L�"�,�9�{��2$6�sI�حЄSZ�h�5L��p
� �AH��1�����m'���h$��ޝ�~J�,.G[��	�F@�4%�}����b�+gobQ�el���V4zm�!=�y����h�}?�.�10�.�	�Z54�݁y�k�����}/��)
��4<�h=Է`nӸW�{|����u�	H�N~��v�kC���r�O��C��0��]�)හ��I��pg���P�A"KۙJY�7C��H���`\����~�/���3�+��RL�a)'r�Ӟh� ��I�;��mȨ"2c�P*�^�7C��Ho��B3�;T������v��㡝�r�O��C��0���t�J0v���I��3Qq�^U�|s.�!�zg�Z�$+�~c(�U���.�O'�W2�����`�f��ϵ���Ԃ�W�o�r�O��C��0��ד�̟a�,��I�U�߷� �9��0-*�&�!�zg�Z�$�H�`}�f���L�B�)�g��I��fP%�SyI�D���i����	x]�������7��Mv�9��a�{�0�!�C��jџ�_�v%�#���{��Hl��f�� ��C���)����Xz��BV�;,J�l�/���D��ܒ�L�}��B���s4y<le��^(hO�Ԏ�G�K���y�\�ʆ�In��t0�'�@ip@{,�����O�Ԏ�G�S]�����<u��w)�S��X3�������Φ�8ưc��!?���5"D7n=������{wÎeT�?�)h�52���,���+�k�8���҆�|n���:�o�E��Y�����rw�O�I� ��ѕ���Ϫ+2��z�W87"�o�9���1�r�O��C��0���df��/w���� �b��j3�w�>��SU��Pa�s��_;%v������J��\���a6�Ͳ
�3�K,��,Iw�)�D���i����	x]�G�Lm=�b�7��Mv�95�KP 4Z,�&�$�kyKџ�_�v%��"3<�Q����AyU��Z��G���Q��ȎC3	^Yt��m�ep����`�����F�*�h�҆�|n���u� �(�ⱃ�!�QD�:mF�'YJ�Й�m���K#Q��-�Q�\M������L���ڰ�]���]�����Uˏ

�2�ո�R@�2r�O��C��0��$�>��w�*��D����Ǳ����w�>��SX`X�B%�r���7ȓC�-`�e�g��!��x���� �"!B�������.�-���
E�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc$��+�{c"G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s���ħƿ�9c:��{~v_z�m%̼�{���_��w���C3�k�����ΈIn'�J�gs�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S�7���I�ri�y�!�3]o��in�m��+�<4��ˌ�ň��h��]�F��������X�f8艢��S��������Ǜ岦�%I^��������D	��U�q��w\F�w�����޳x G����^������f�j�7ص��s�r�X�<\�%Ah�%4
>��f���T,}��I�d�|��6m�������0|]<w:��b9�����9B7��QeRx�eg�� �vBX�y�`4Zp��/����l0��F��jY_���P[���F#gŮ"ë��}�qJ��I�s�(�ߜ1��b9�����9B7��QW��2�+�HUv�׿e_=����Y.�J�4�e�(�4q���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3f�X0����ߠ�p���R*��7��As?~�F߳��id֠���ry��_�J�c_�;��㹍g����Q�<��׳�x�g�Ŋ�VNy���2���,2�]���/1(�"Hp�,��o��9D+`uώ� ��C���!�`�(i3x�]�V��!�`�(i3��d҃!�����4X%�X]q������>�qxm�N���֜x3ֺ:v~E�)d,�ː�rn�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�-�W��������Uo���<�K�iJ�[�u�:�z�4���D+`uώ�Q��s,�~TM�e�w�G������i����D	��U�q��w\F�����n [�ܺa&����1�9��`�ox!�Q�W���`~�ߪ �)	�8V�@Uo�\/QD�v�l�Ū�TD�����u*K6HY_���P[��I��};y	�Y��{?a� ~>>ը܅%Gbx�]�V��!�`�(i3�I��h��	�Y���1��� �U��֜��3JHn��z��x�f7﹏3�{z�k�/���i� � �	{��Y��
�iC�E����F��j��\w��0]��0�&�ͭ�zT�/�k��j��\w��0]0��l!���?�{�T�	yhPGl݀K�6[��u�a�*��R4��-��%Mό���.�U����ޚ�w��0%����-��%M�rs�i���`�M�	=̞��>�B^`ٌ��x�[5��Z�8���/�l|�*"k���(ӈ���m�r����0C��؆Q>�[G�-X�@�^��1�0M�Ŷ�8k�(�y���]���>����C�/$�ߺ��]Z���W��dI��w��,>����C�)��7��Y(�׿�߼�E��]���>����C�8aPe��׿�߼�E��]���>����C�U�0��IuAw�8�}?��]���c�A�L'��~�2�?؟�r�`U���6�˝Sz��E�4.@��/�G��x�8���/�I<��fҹ�\�<�dQ	���qk�ZV"���:��#tC������s������n`ۺ������Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�$:v��`E�EYZ/�h�@�o��I�?g�f���\X�<����8��U�/?��qᾪ���>��9���$1mp�m~|�քY��:�襈P���y���JHn��z�qz��u(��@����gGɑ1tc5+�o���B���+�J��P/;D����L�E�$����Y�Q w�)/�L�He�-�c,!3�?4���R;7s�9���o�jƓ�[����ըi:�HCaIMl��*�>^&9@^7&ģM�I,�D�y:#9�]�B���' ��Cҷ��ecx�S�����S8���IO,���������9b�S� 7�v�ԯ��Q[R�7����n9�O�M:R	�d2}�#�l�1����?��/��q�&��DP֞ �+`����Uзq8�Ј'���Xw���,D�������z�
1���;�n`5�fK�\w��0]b!��uፀ>1J��� ��j'�S�]�!��	Ǹ�y85�B���0�1���U���&\VI`,'������݃�Q[R�7�>D��e2���HF3}�
�?��&��>�!�`�(i3�d�٣���N N�S��30���,"�x|ٲ�зq8�Ј'���Xw���,DH�v����ܕz&�8�n`5�fK��0z�cUL���.�1�3�8���/����,D�x ��s��q���nm�n`5�fK�\w��0]b!��u�s�Uo���]H/��d��]�!����w�Հ��}�a��>�A�IS��#�$�~�M�q���U��@����gG5m�E��P����z�7s�9���o>��l%i�-�n~�x��͘D5���E����FZ鎬������_�,�����?�!�`�(i3%Ah�%4
>*"v%)��2�����B^`ٌ���C,�V3a苯ܪ�\,�R���N�����5\��{��G�y��s��w�q7RSJ�J�婎^���y��������z-t"wdC���O���߼
�d,ܕ�21��@ ��#P�^#9�<�H`�ɕ�����a�"�fE~�c���zU�[�?��J�8�+�
�c�~�Z�>)��"�,�>E��'����E9���R�փ(R��(��$��Xo�dI��������D	��U<[@�b�����T�����my$�N�R( y����Qs9�ڄtm5��1b�N}�m��{ȶ�k�7,��n`5�fK��0z�cUL(����m���omw"$/��/�I����g��v�|[��N}�m��{��Bj�F�K}�^<o}?�0z�cUL(���O�!@�O���{��~�26��\]b�"x�7�ܥ��2��[����J��4W��C ��b�FP&�%k�����d�٣��c�A�L'�}g6��g�s��hq`�(&�L��\}{��귡<���Ŝ�	��"���>(�6k�4d�>��m����[L@3v'{w#/ B���#�cQ�H}�c��T��a �5�6#-��g� h�ҩ��'�PN��dN�<@Iv����-�T��:5A��p��jVѭ@���M$��v�@����b�z'hۉ)/I�wz�i7mŀ�\�gb�r��>!�`�(i3�E�F͏G�Ro��IS���m�������F��O��|#HK��55���uMA&�:'���Xwd�n]N�F��z����@��v{�G`,9�H�WU烸*={���	�|����؟O��Оp��pZ����C�c������{[� ��ǐ�EV/^W�"�!�x=�FZ�څ�?k��K��ʁ���Mյ6�4fO6�e	Ղ�I8�y\��S��z�m�QA�Q* !�`�(i3U /숇�3���U��-�;S5b	��T�.���NM�����6�������)��U젩`#FW8�	��y�aC;�}Dq�f�G�&ց�*欄@���tn���}���S.�3�����s;nI�!�`�(i3pı��0�����G�VƄZ��3��w��\�W݉���H�,��ݓ�W����Y����|�4�0 L?ஹ�%�Ԟw��c:�ݚ�Н�(*�O�qF�Oz���[}�N�`2���K���Ѧ=84u!�`�(i3"�+yz�T��&~e�e��E{��h��L<�c����|e"ʁ���Mյ��5e���A	Ղ�I8�y\��S��z�N�G�,�!�`�(i3U /숇�F�>0�)-�;S5b	��T�.�ӟOi���6���X���l���U젩`#FW8�	����&8nm��}Dq�f�G�&ց�*�֖�&G�n���}���S.�3����t�ė�!�`�(i3pı��0�����g��dބZ��3��w��\�W�����1��ݓ�W����P���4�0 L?ஹ�%��A��Umh�ݚ�Н�(*�O�q�b|l�H�<�[}�N�`2���K��&RP��٥�!�`�(i3,�n�a�4Q�&~e�e��E{��he�<�ڠz���|e"ʁ���Mյ�$0B2s�	Ղ�I8�y\��S��z�</�#���!�`�(i3���'��@�my$�N�-�;S5b	��T�.�"ث6z[fĉ>99��|��3�fĉ>99��R�V�"�0�[��p#ِ.�d^�ϓ�������`��5ߧE4��O�{��&�~�������Z�{/J�ڙ�$�e�D��cEp	���>P�2-i_q?�y�I����h <{>w�\[��l�,U�Nj�N�R�7ʌ�J1����?��X�K{�(ms��/�u���4���O�>�k}�r�����Uh1�;��|B6ϔO��)E2�DZ��L�T�t���O	��c��B}�4��d��D24N<I8����\.W^�V]��}���_j�Nh�EC��Q^�MY:�~��;�,w�R���y>��yСQK:2i������ÂY�`�!1��L��Nz��U��)��}q�k����:���
�XDt����VjԿvU�E����Fxy0�u��¤M�[�g��DW��ԅ1Qr��[��l_ ��b�FP&p�]f�"v!�`�(i3���#] ��2N��n��ޜfbyQ���4���`��V�^3C���_����$�Qu�R�47��vL n9-�N�W�E<HӍ��`���oN}�m��{zh��ʊw!�`�(i3���D	��U�SҤJ"�^};�ۑְ���
���}�D24N<I8����\.WX3�������Uh1�yO�E���%�;���EWr�!�����"�,�>E���Ԗ/�����IO,��������;�¬pX��g��U-�e�,���6+� ��b�FP&g�P7�#�!�`�(i3jݭ�F����μ<�e<�.��|ȃ��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ�F�А]��
�M����d��-��!g��J�s��z�
1���;�����u��r��f���Ն� ��%�D�v�l�Ū�TD���7��y%%9���.:��Q?M8�f2!�`�(i3����0�������ߺ��8�ۦ�P�X��P�������pC-��h�>
A��%�.MB^Ms\HqWU���>
A��%�������}� h�ҩ�!�`�(i3�����4��aP�T
�k�:�l.��L�1p/-��N�]|-��n�_*�!�`�(i3a3@��[/�L��O��p���[`�K��}Dq�f�՝� s�#�BB�k���1��� �U��֜��3Vr�O���J�\���=-�aT���ǧ��b�@Ñf�
����J;���[�uV?��?s�̵�7�!~u��r��!�`�(i3�g��2����͆���_�=[���:�HCaIMl�T��G,���ݚ�Н���6������S>�35|F#�Y
�T�r�5�!�`�(i3\OW�:�ݎ�T��ߌ.�� 낢Rb��Y�WA���V?� h�ҩ�!�`�(i3;Ε^����#��ߨ{���Γ8��������t����>PQ%cp��g�H���~��!�`�(i3���F1������$��;Ε^���3$�J�5'!�`�(i3�߆�p�hؕ�V�&�>
A��%��䓴�l�(�)	�8VڂK�ykv!�`�(i3�a�}�$�
Cj�R[z�(�� '�i�*ڶ�UKs,��L�1p/-��N�]|-��n�_*�!�`�(i3a3@��[/�L��O��p�h].K��e)�W�=�k��:5A��p
�:qEp�;�P�t�5!�`�(i3<���K<�Vq�|`kK��I����<����1tSjv�!�`�(i3���F1��kټ�b�	�RCJ�����@�ĵm�ݚ�Н��Ra])n#���r����!�`�(i3ml@*���'�ɳ��!�`�(i3ؘ%��i��"X�8�`Ut��\��?��a-�a��@�7�!�`�(i3��6������S>��LH`y
�{?a� ~>�}l�c���}Dq�f�!�`�(i3�5ߧE4��!�`�(i3HN��R��bP�63Z�t���%>�rG40�RS���$
�)!�`�(i3��u*��N���{��c����'�u�
�B� �b��!�`�(i3���F1��kټ�b�	�RCJ�����@�ĵm�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx4��<��^4�1�[;#��Hۭ֯���,���#�e���gmJ/�� ��b�FP&Qi�d��2c<���z�wnB�K���X��b ��b�FP&
�E�6�g�Y��]����Ż?�N��+x�r�s�*�I�x�?� �"5� �St-p���|�d�G}%����3f~(����[��l�,��ȻK! ��5%q���f�e�M?��yЈa�}�$�ϔjZK��#��_�?�tT�_�X�p�cȓM�Me���F���A׏23��;e���`�{�P�1|�����^d9	��l�vM�=�~�Ԣ��%��J1C����B�+ty8�:����G� �X>���\4T۪�؉_�'���~� ��S6~4@ڲ�.j�G� �X>���\4T۪��N��Ĺ�+�t2�֯���,��e_c�?D�8���������+�t2�֯���,��e_cƍ2���l�\���F�`y]�ś�'��x�`El�H�RtV�^5�����}Y|�l<�K���U���t�襈P���y���*A&-�Ri!�`�(i3__�n3	r�(�L �Gȇj�Ï��	�.���~!�`�(i3fF�5.]����}Dq�f���Ě�����}Dq�f��5ߧE4����R��%4��"S�F�KD�Vr[/}>5��0$r�t�}i'{w#/ B(it��0���G� �X>���\4T۪��N��Į� л��o�t��z�
1���;n��뾦�<�6�Q=1���~��+�t2�֯���,��e_c�?D�8�鈥�J�a��.Vȼs����R��%4��"S�F�KD�Vr[/}>5��0$r�t�}i�;�P�t�5�׹���C���N���7�|A��O��� ���Ī#q�0B�6�o8:4�I���c�90Mj�dL�{y����i�q,?5qTdJ�{�yü(5D'����"sS<GYqcHTX�';��#j��=����t��¤�<TC*���H�e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ� ���Aؠe�:
1���Ư����z���!*��*8�N�Cٺ��#o�]�ʄ�ݟ�e��Z<��A!��-����!�`�(i3�>1J���3�Z�Dg
�Pђ�-�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�B���ؐ1 qM�[��Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���jA�)�H*�^ݙ.�����߈j�N�p�`��g���rz�rX.桸���0�G�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT����ge�Ip�K\�0�U��)���yk;��2N��n��bcb�q�\�K���&���\�v�g�W�I吱 �']g�׺�&\VI`,;dE`r4�����+�^n=\f�5>�y_ G[[���n�".�\���F�`y6\�4�@�� �-j�1tSjv�(܆�NGV��}��6�8�-Zy?X���a��ݚ�Н�}���yb���}�@���_rS�b�8Z�AԢ�a\�2}$#h6������t�_�֖�߾����k$ �����i��J����[���G�����Gܘ���a$f��_Ub�F�S�1 �s`<ܧ��M/����A��'�ɳ��!�`�(i3�l���dW�"/��@��s)9l�R��0����J�Zj�����E|��d��R�^^����s�Uo���,ܓh�,�[��hg׸�� �?Ct���g[��p����y��j�ɋzò�W-�����A�M�Kh�𱍞3ƥ��_�_P�yV��>���~3B��%:�d��R�^^����s�Uo���03�� <I[��hg׸�� �?Ct���g[��p����y��j�ɋzò�W-����Uf(sh�Ӏ𱍞3ƥ��_�_P�yV��>���~3B��%:�d��R�^^������U�R^p���P#d��:Etj�/��@����	X%+�=�x�N�M��*�8��S�҇�8�\���l'��GHS{�tץ���q�H��{���U���C���C�7�/�)h���Я Y;�Uʮ�V(YhV|_��{���s�y��j��k$>"A��⸱n�����?��#b�.]����q놕
�C��յ���fh����p���3�eO��W���[��l_�5ߧE4��fĉ>99�� Ӗ�t$�)�vxy_ G[[��K�ί	�����)W�{n{�V,���?6ֵV�-�N��8�$W+͝�!������t�T��?E-h���U���e��_	�Ƽ��S�J\72�d�6?�;D�Vh2G�,��R(�U���e��d9=���u��r��bƑ��M2B�FxUƍ2���l�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l��L���;��81����O=�W��u]9�#�I��-����!�`�(i3�����o���8.��휯}Dq�f���Ě�����}Dq�f�}I�6���N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s�)��7��Y( z�P��1tSjv�
�:qEp͘D5���q9+t�}�ݚ�Н����F��O��ݚ�Н��5ߧE4��HN��R���ء�I��߸��S�Ȍj�����)�_�D�s�Ư�ճ�%6�E~K_���k���2 �4"�ed9��+����$��r����!�`�(i3!��vΣ�wR��T��<l{�]&"("��ͼ��!�`�(i3!�`�(i3!�`�(i3�����!�`�(i3!�`�(i3���۸Y-�D�D��b���|�Ȝ�ɵ-�C��7�8)���M����z��� y��,'{w#/ B!�`�(i3�#N������8(|8d�+Y�6R��M�,!hޖ�A$�P��O�@יߌ��omq�:Fa�7��Ɨy�"c�t��t9������"sS<GYqcHTX�';��#jPM�^-qXi�G�y��)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�B� �b���H����o�γ�ha��o���H�RtV�^}I�6���N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s�)��7��Y( z�P��1tSjv�%?gV��UXi�G�y��״$(�>g�
�:qEp�;�P�t�5����l�� ��5%q���f�e�x��w����֯���,mk��L���R��3���Q:��?��a��o���H�RtV�^J>zߋ��>ַ�����ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}���$�uG�N6-	����+utM��楱�o��_�Rv�䩲$����E)e|A��`���φ��<�6��&��>��7�癆cgR������������ h�ҩ���v[2�'�^��������@|����^a�nu4Bޗ��jw�	���|#HK������ �'����u��r����#�a�Ą�ԬQ����5��t�	���QC�꠼*d�m�d��-��!g��J�s��03�� <I�����&G!�`�(i3��v[2�'�^�����ݚ�Н����F��O��ݚ�Н��ȟ�P~
��N�Cٺ��#o�]�ʄ��.�L��w)��
=b~*��s�)��7��Y(L��'p����-����!�`�(i3�N�*��	@%��v��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�MR˿�lw&�;}it�<��#b�8�@�0p(�OZ�'6��o��r�75L�`���6���o{b�ʐ�v��7�tɱ>�����U��)���Y;e�iK-pm!9�>��n4s1�U��B��-���忔8��;	ȕ?�7�癆cgR������������ h�ҩ�`&c�'N�j��O|���/��kOT*qA����6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i3����,����0�|섃Va�ir=5.B����1F#�֞q�<nD��.ama�`m��-����!�`�(i3s�Uo���ַ������?D�8��HN��R��bP�63Z�tL��/\�߿�wW���Z<��A!��-����!�`�(i3s�Uo���ַ�����ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}ĚȜ��Y���ۉ��K�A�a�ܥ��(J]֞��_�TYh�p��_����3Y����P-r�uh����s�Uo���P�<�^�s�IX0F�MV�ҁGG�K�BN
\�N}�m��{|�v�����G4aL��zL͊�q��D2<�4j��`���φ��<�6�`&c�'N�j8D�r^�Hd���"sS<GYqcHTX�';��#j���*y}e�����ӽC�H�CW8���[{/;k+Q�h'�Ȝx�5W ��̫(� h�ҩ�:
��x�{�\��N�Ś�-��������l�鑴HH��"�̙	,N��>�s�,�H��-����!�`�(i3�GI�\�0�c��v�'�i�*ڶ�UKs,��#��I2�8� S������v�9�ʉRa])n#���r����H�����?�@,��V��J����(�ߜ1���}Dq�f�fĉ>99��A0ok��!�`�(i3����,����0�|섃Va�ir[��l�,t���H[W?ى^���!�`�(i3=|u�0�#1��Z<��A!G�j�:S�Lm�<o�̽���z������ևA1F#�֞q?c��qg���N�T?w�;�,��1tSjv�V�Ո�����������4Yz����|e"$f��_Ub�F�S�1 �6�>�@�	�ō܈��V z�P��1tSjv�V�Ո������ӽC�H�CW���|e"$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vx�m`���ZXH�7wS��h\K�5~�Uʮ�V(YZ��*x���`�p�*X"���փ�ӇciW"��,����ɮ��"�*���"�k�&��3C��I�(�w}�tM��楱�o��_�Rv�䩲$����#��i��~�26��\;��B�lXm��G��*IÙ=�HV%~YqsوiI9�o«IX0F�M�Uʮ�V(Y��a��R�7�癆cgR������������ h�ҩ���U�R^p���P#%��v�ڹ߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#��"����G��Hb� h�ҩ�.%ĩ.u:�J��I�s�(�ߜ1���iB��H�RtV�^U����ޚ�W�o]��e���Γ8�dKa�����Q؃�L��r|����$J�-��^�Ra])n#���r����U����ޚ�W�o]��e�����<+yj��x!�`�(i3�5ߧE4��!�`�(i3[�5���78�íN=]b~*��s�/$�ߺ��]���޵.�ۃVa�ir���ևA�d��-��!��:28�|��Ǎ��I4k05B��-����!�`�(i3�Uʮ�V(Y�t���1�g״$(�>g�
�:qEp�;�P�t�5����l��b���G�ɥ�|�Ȝ���'����u��r��a�}�$�᢯��0����$�a/��kOTfĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�
r�	O)�A�IS��,�د$��ѩw���]�T���A�P_,�W���&�\D��D1��n����ݢ������쒃\&��Ϻ��S����=�Uʮ�V(Y�$��fG�a���t�T��?E-h���U���e��>�2���u�#��nt��F�z�8#�b9���:&�>��s��n4s1�U��B��-
r�	O)�A�IS���=Djw�9�xjzӝ���w3��׍�&�U��f��a�}�$�᢯��0���O|���/��kOT*qA����6\�4�@�� �-j�1tSjv��
�t��T&��ۥ`�M?��y�!�`�(i3��T����4.�ԫ�0�	A���-/a8!�`�(i3��N�T?w*��D�x���Q����.��$����zܳX��Hpt����}Dq�f������!�`�(i3��N�T?w��OZ|��������Y�I��fĉ>99��A0ok���H�������+1�;�.��1��!*��*8��!�qgy�`��vN	���QC�ڎC�?��(4G��>����#��<1tSjv�X�o|3bK����ښܔ??�"��ӌ�r���%>�rGO�D mWN;�jmT�#��U�R�ܬ�mоG��Hb� h�ҩ���೹�C�A�IS��ַ�����ƍ2���l�HN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}����L�yEB~�S;�����*��>zƑ�i^�U��)���Y;e�iK-pm!9�>ֱ�q�����ѧv;�?�@,��VJHn��z��r9�3d�G}%����3f�m����2G�,��R(�U���e��d9=���u��r��u�st����'�PD�����g�Z��3��a���!@�f")u��r��$XR�QܛOcOZail������&G����l�鑴HH��"�̙	,N��>�s�,�H��-����!�`�(i3}���yb���}�@���_rS�b�8Z�AԢ�a\�2}$#h6������t�_��ݚ�Н���jVѭ@!�`�(i3}���yb��-H��.�����o�����[��l_HN��R��bP�63Z�t��#�a�Ą�ԬQ����5��t�	���QC�꠼*d�m�'����u��r��;�jmT�#>�{>�Ч܂�F�z�8#�-�ྜྷ��H�RtV�^�"�чE4�]�p� �!�`�(i3�����!�`�(i39O�m96�o9i�!>������fĉ>99��A0ok�ª���l��x��V��y$�Rt���X�R��3����'��8k��.ͥ�H�RtV�^�"�чE4�]�p� �!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f�)�{6�U�����F��O�}�	76�&�� Ӗ�t$�)�vxyk���]{6�ǌ�lA�>P�2-i_m�;Y'�V!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��F