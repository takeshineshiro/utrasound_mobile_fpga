��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag������T�h��~�a.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I��7��_�L_H��Y씤`��p�eh���w1�I�?g�f���\X�<����8��U��Ĭ���^W��C*z�w4G�� ��d�n}K-J��K��z������3�z�ω���D���+��O����F72��{L�8br�.�/�d�������4�;���u�$|�>I��4�Y�YrT�#.�Ő�|��h����jǎX������n�q���xP��t䗒�|'r�tI����j�6ˊA뫕p)1 T�V	�tL��	�<�A�}Q@���rahH.�J#B&ljW�n���8�U��]>��D�,�Hc�.[K��m�X�'b�mh�@� �ʁ��+��| '�]f+P����?#�+Z�q�PO4V6��2el�h�зb� ���@��;4�zu%��HwF�E0�G����/�t6~z֯{�sg*����wx0�<����ʉ�����0!B�6��[���(/�j��⫰(�[6L�}�2��N��4�ޜfb��h"����P�Lư��I���[��@	&�~��F���	x]�G�Lm=�b�7��Mv�9COŔ}B�+t�%A:�	8�:r&@�@S����a��F^Ie̞fG�a��un��H��eu��w)�S��X3���7��Mv�9�'d�
S�u�
˞�|�8�:r&@1�+Q�<�pQ��G�7�N���D<����d�kⲬ��;�Ӏ�I3��(���\�4�s��{��]Q�TT	q��$|���Xd���>ӧ��~�MUs sg2^�L�n,��J���h��W���4IQmX��d��9")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�1��8�h�� ����f�#�eM����c���o�����0��D��L���_�L�Ȳ�V�溜��D�,�H�R$�� gs����'v�]wɭ�7��r�=!�`�(i3N�By3��<�]�!����M[��Ǣ)�k�4�U!�`�(i3�����5	���]����,�JL����?D�8��R�����!�`�(i3�����5	���]���>����CΌh��eZ!�`�(i3Y%T��BPe.��xu	�>��l%i�-�5`z��s�Ƀ�?PA�':E����j���0z�cUL�I��6���T�\ ��:E��]��8S�n�(�a�x�f7﹏N�By3��<�]�!����M[��Ǣ�K�&�a���i|�l5R�����5	���]���>����CηxmQ,ۘS!�`�(i3Y%T��BPe.��xu	�>��l%i�-��E/��FH=Y��@�E����F7G#+��\w��0]�o�t��F�e{iʖ.	��A���TD��ό���.Ӂ��̰�!i�q8�2t�ݡ��1����(�
t��Y�{'%s2�ew�a(􆿳����^���(R\֎u�,��7-�)�V�3j@IE�U��>��l%i�-�jo�'q�!�`�(i3�E����F7G#+����w�V�"�"��FX1�������Pc��q�Pe:[e��m�D��L���_�L�Ȳ�V�溜��D�,�H�
~�d�9��0�S�&����B	��Hk3L~΄gO�3ׄ��,�&�{C����^�1�:�Ω�s8�R�	�}�����`h�ag������T3ų�̿}�
�?�	�%��6�1�#��d_�n`5�fK��@5���<ZJ�hEc�>�T��u��!�`�(i3��Q]� _ό���.�}�
�?���\���S)��p�:��n`5�fK�\w��0]b!��u��K�&�a�PB����A7s�9���o>��l%i�-5�e`��9PB����A!�`�(i3�d�٣��&����L�s��t#�z��?e!�D��u�(nmm�`n�m�W��"jm�v1FL��L5ӥ���98�
x�?!�`�(i3�E����F�5F:	�����A���Ws�N"T8��$��<WNPB����AlC��ۺ_~5�Ǫ��3 "M�yVW����n,��Jdw��D����úAV�!s��V����3ɂ�δs��t#�z��?e!�*S�jH�}L5ӥ���-���f����Oo;����V������D	��Ux8��捽L5ӥ���-���f����Oo;�lK9��F�C��l"�u���FR6niܒ������b���ν���1��v��OD��КK���4|��!�C`V�-(�e<�ߢěf%װ$��_�W���t�U���e�AqeGfB������kO�%5�����Wo���˃�e��������p1��`p�~(�M��1�, ��XJc����Y\������*��� S�n�(�aĆt$�(�\���>�(��G rgA�iK�D�b=��p�:�F!��D�����k$ !�`�(i3!�`�(i3����_Bn��akF�e{iʖ.^R���	���������d�O������lĆt$�(�\���>�(��G rgAS�n�(�a���3E��ާ�����ݚ�Н�!�`�(i3�y��j��k�BT	��.�8c�D?n�D��u�(n�%����`��g���4�@	�u�azG�_h��]߱��qC�G����]'\gWg��	�Z�kfcj��r���iI9�o«IX0F�M�ȏ֦�"�\���F�`y������T�8k��.ͥ�H�RtV�^g�G��0RR6��-z��ic)�̩�?D�8��%t̓�@�O����&{�A���Je�"��ӌ�r�i+��_1�f���!�`�(i3n��뾦���l�^!�K�g;�UA�qIp��K����c
=^Lma��Ck+Q�h'�Ȝx�5W ��̫(� h�ҩΪ�\���S)��p�:��I����~ug�G��0����[j�%t̓�@�O����&{�A���Je�(R\֎u�%s����K7�wtMMRR6��-z!�`�(i3s��m�Eq�ȠȎ�8�ݑ���&�d���%O�	^���y�%5�����8��"�7�y�b�G2$f��_Ub���uQL+��φ��<�6��]߱��q�� f�0vA#&��Q-�b�+�