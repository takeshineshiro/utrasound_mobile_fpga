��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVD�6�����;��sD���L��+�Uz�QL�]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUP���*+�[��������-�7�5��;��sD���L��+�Uz�QL�]��;�I�����)O��Ξ4�"�\�� ���K�O�{����ۤ�9is)V��㝒c\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<���-ZW�k%u�e<��⪘����t�켻�S���c,� � U�rN�3��m-�@xI+r�� 0�D�A�f�mX��)D�b@�WVJ{4ȕ�c������j����t�5����`K0�Rճn���8)K�h}�Z�z���	|H��z[�wf)�y'��BS��TC�w���0�O!.�ޭb��G����a�����(V�>!�/�7��u���nEA�����5O|H�!���Ȗ��h�}D�8����TT	q��$a4�����i�p&�K��~�MUs �c㚂��T
u�/%�ĩ8��[��`�3r�O��C��0��`�R&.1����_0e�v�h�u���;��.~�Gj'$�o��'j���j�r��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���4*�7\��4�/�I����D;���N��j��D���s���ħƿ�9c�1��8�h7H�u�ÍeRuw�C?3d/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_E$ô&y�#�̔"v��ƒ)?˳ea�8����]��
��rE���ƪϤ�Yk"1/Y#_Wӆ�q�©���H��JnXe�+�Uz�QL�W*g;XcdA!���oV�>!�/�7��u���nEA�R0��Mfp�m~|��b��}�����ތ�1��\�v�a�fj �.2��m �A?��V �-�>&�&i�Ln��S�WT�����NuG�פ���Ћ�l�T/��=��K�Q��T��zL͊�q��|�&�'�2��m �A?p\匔'�?�R��nDK�e�PV���\�v�T?�7G|`�$��Xo�ab�Afz>��v�8:v�`M&3���\�v���GAџV�$��Xo���{�3�P���ġ��,Ln��S�W0�T��:hΕ���iv��-�2��%�/��Z>L��n8���ٳ��溂�U~܎VV��5����`Kְ�4'N5wĒ����H���o��qo�:��7��k'�w�������O�Y�I�4];ˍH���Vch�,�?��V\����iW5լ,� �x�]�V��w�7qyX�񙗡��\���,�?��V�Ћ�l�T�r�&U���0��PWLn��S�WT�����NhΕ���iv��Y���������u��rW�#�ڊ<?@��[	J��;ѮK�M>�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�V&����5����`KI�J��#Kl�Y�7#�xI���|�r�HzL͊�q��C.W26K�~��^̽1��H����8�A)�V��/7��k'�w�QP��=Ch<Q��T3�2��%���Ặ��Ϊ�Q� ~��7��k'�w�_�s���H{װ?�p���H�MPq6.JHn��z���G7�����Q�bI��'�����7���{r�����ތ�1��\�v��D�����H�g	�Ϊ�/-T)x�?{���x.�Knq�ɿo|��g+��tI�F�;���N�+��o�U�C�u)�6�Օ��qv��3�.�J�}�|�݌��r��VYW\-@��F~*7���&�_0M�/�s���'n�^0o<H�-��*p�m~|����� �ܰ�a\Y����)���8҉g�kG�#JHn��z���z�O҈��n>�ϸ��Ћ�l�T�I4��欱���j���Ln��S�W�.�p�2�zy��#Q�ܣ��J5$��&l����~��=�����A���ۖ�92���nQ�rVe�Y�gtH�m���E�Y�!|�α+�5����`K��M����A�m�(�^[_�e��IÙ=�H��Ӿz�Vzy�g���+;��7�"� ӫ/��mk�79�����Ψ��F$��O�&��n��l���a��|��Z�ٵT9L�sJ+�e%ސc�g;�C�2�8�aq��@�)d�8��;���N�i���
ON���:�hΕ���iv����	�vI0���ԏ�.fOe	Ln��S�W�כJϾ�ig()��ikp���H���F�-�Xu��<om�����H17��k'�w�]a��1qh_�n�To�[r��}k:���3xļ�\�v�����/٨7��k'�w���j����rx�y�Zgl�?Z����JHn��z��e���0�m��6�~�N������ߟ�|Ń�8�2����z2/PN�ǁ�f�T٬�����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�)��\_��f�Nd+l�Yҽ֗�ҹ�>a��G��x�&[�ͧ�?Y;�L���9�D_�3���U_�+X�܄�֝���b�Bϱ�����7���{r��'6���;8=�g��U-�eI\�53�f؀qjZ�`�|��K�z{�x���;�L���9�D_�3���U_�+X�܄�֝���b�Bϱ�����7���{r��I`1R�J�On`�(=�T�\ ���( ���S��%'�q�5D�=�Tmc^���Ф�!~;��i�̥%�CvK���9u$d9�w�"�Hߢ�<�ȧ�Z�'6���;8=�g��U-�eI\�53�f؀qjZ���A3�(N��㎏qló��|�����V��ߝD9�{��灊�O�i���Z鎬�������(���`$�P.eE�ƃ
ᾆ�x�T�\ ��D9������z�C�f�����/�|��(`��ү/�O'�=�1#��Z�����XP��ȇ3
�v�v-}�	mp��.
����.ᬵy�����b��Ep�m~|���\��j��<%�a���k�79�����\�v�ʋ Z4.���A���ۖ�r����2E,�J�|Rf�� �hΕ���iv,�v����;^�6#9�H�MPq6.JHn��z��p�Sg�3 ���t��f���j���M�I�h�
MQ9�F�hΕ���iv,�v���&��A��.D�3�%x��GD@�F��q���i��6	�4bp�V3���[�ͧ�?Y;�L���9�D_�3���U_�+X�܄�֝���b�Bϱ��R<�����á�~O��L;Л��|#9������/��&����H���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8����ٺ?��+���LQ���"X��[��Q[R�7��)��� "��O�9��+�pDk�W+`�x�o���{��&�e�5
��ָM�n��ҹ'-����-���p�m~|�֯f��[9u�Լ*�ꄐ����3mzx_�����K�J�ɤ�ud��d������yZ�����~~W/�~f�E�L�l'�l�p��i��C��O/OJB�D|�I��'�HaU$kX��a\Y���1#��Z�����XP�����w�K�1c+������U��+�X�{�5\-pD9������$��Xo��GR��)~s�����j�|��IÙ=�Hw¹��<d��A^J�po4��;�vL?���3Sރ�+�c��7��k'�w���j����r���*j�B3g�����zL͊�q���Z����p��R�}vJ^k��Nx�^����X:L_ؚwP�+mw�J�^�5�a=��τ�>��I��ɬ�[��ZݜC��Q7#�6`h�5,Wl�/�O'�=�U��I�v��s�h�
!7<���������	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�/ #O�)Ĉ��r�]@P�B��X��8���/������Y���e����0���h�����zE�s��3���'ɮ^�T
���[B.�OY�]�$d�I�v�w8FF��!!@��B�֙D$����m�p��%��Fc�Q4R�q��I�X�fL�G�Ȃ�8*Y�A�Tl�L��M�,���	N^�U���%Z�*�p�m~|��8yL2�����ތ�1��\�vŶ�T���Ĉ��r�]@s��I�λT�v��1�; ?��������n �9� �Y[-t"wdCu�!uqE&^���:r:�hDP0d�� ���跠Ћ�l�T�(��ԋT���S���'n�^0o4��t-s�e�J�Pn\���k�(��z�u��hr�2����<m�M�u���Ϙr�P}؛'(� B^�.�ߘ�)�I0M�/�s���'n�^0oPpkiq�o�H�MPq6.���fa���ӵ#yӛp�Tr�j.`#2��%07��k'�w���j����r2��������������JHn��z�>�ack���A�;�֋`N(��/沄�J��CK]���.�#�0!S�,��ш�A3�(N��㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���_U)�<�&#�+���LQ���"X��[��Q[R�7�ͭ����f����0+W���F�^��NP�b9������U.6��̞��>�����Dɵ�p�AJ�e�$�,W��+�Ds�`��=i���Կ,��_Vl�A.;��L�O����K��p�m~|����U0����d5�:�w�+���LQ��b9�����:�{��ߘ�)�I�3�"��+W���F�^��NPz5��*t����eR��C�`�/�t���|�r�HzL͊�q��!7�dߎ����d5�:�w�+���LQ��2���O�w(��ES���v�8:����P'F2��m �A?�����zPuZ�v|��3�%x��GD@�F��q��W��Y��%���It�Ɍ+8�3��$<�Q�R�j�`��2�.�05k
��F�2�q#O��*V<�ɔ�u�I1|��q�����]��aT��0F��� }}�@ de\�x�ҷ�������?ןuɬc��WN4�CL_܆$
�L�)
`[~&�x�$��Xo��_��f$����ތ�1��\�v�h}{���wk����׃�Q�.�I��'�fÁ��/�ɵ��!d�#�ڊ<?@Pʶ=���u� ˂c�Q!G�bk����{UGICe�;����J>п�p=	�˳͠m�xW��9u$d9�cx�S����jƓ�[�$��Xo��� ���Lk�Bgt�#P4];ˍH��M��=�&&ĕ^$&�	�s�{ܰ��G�&�tc��P9P��`�.�D���J7"z�T���p�����õ���:�v���p�n5�<�a�փ���@��O���Қp%�&zΙ�[؆��Sw��9�Vj��84lZ�Y���W��v���s�=��hӕ+G�7�mEi$?��ז��n���f���n���|�(#FECJ���wb�S��V��\����X�N���{儫y����^/�?��H������~��mEx���w�s�v��؄aX܇5����`K-�U�a�&9F`}Ĉ��E����Fe͉�Xk����0������Vϓ�;Zr�î�DԮs����Juq���L���E�H�^�A��5	��������8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��Ź��Kh�����6�(U�6��f`f���b'n�nh�l��w6g�D��l�8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3����e��u��/">Q���eټ}B*%�~��/��l���&�	ݹ���n :(a��2����PD��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��7O.�p���_�e�T����NJ��"t��̳�(<n�`1sZ&(g�[�x�w����N���0�����õ��ޒ[�ɓ��Т+�m�����ܧ@��O���Қp%�&zΙ�[��$���{�����5_����wA�b�V�}؊Wo���>���Ч�گ�$e��'IbA-!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3I��-P�gC+�?8����?rɼS��5ų�_{yL� ö�M+�~��3�-޿I-!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3w��~�:wR��k�ݝO��6�q���ɨ�Y#���1,F�*'&�� 9�q����s����Cׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3c^���d�L���x�cz��lш�R�+�݌�[�y�m�&���i�9l6�·V��J�<'���l�p�m~|��y�= �t�����$^�Vn+G!D��Ψ��F$��O�&�鱔�]�,I��K�D��2e�6��ѝ�9��&n��������QK�wux/.7��k'�w�4�(QG���wa	dx	���S�?_.Q�q�v���{UGIC�ҡ�֔���_c�}v��7
��=�,�I��p�m~|��y�= �t�����$^�,��!Z㘢��Ψ��F$��O�&�鱔�]�,I��K�D��2e�6��ѝ�9��&n��������QK�wux/.7��k'�w�4�(QG���wa	dx	�N-��	е�Q�q�v���{UGIC�ҡ�֔���_c�}v��7
��=�,�I��p�m~|��y�= �t�����$^�BP��ٙD��Ψ��F$��O�&�鱔�]�,I��K�D��2e�6��ѝ�9��&n��������QK�wux/.7��k'�w�����ƆMs�ZoZ.���[;Y���4]�k�1 �O�ox�'g8�(P����o��?#�|��l�dǭ���
O��'��*>S�	�:�F��+'�sȸ�"rR!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3"�(��t-(a1o�j�z�a:��N��ᷠ��/zE1�4TZ A�����8R'�C!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�	]}NL���g����|�Ԏ�JJ6��r�&���'#�*p.���l���zo��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���;#����s��8�R���G�E�.\�����zG�7�mEi$���0w���_�����������t:.0(��6��e͉�Xk����0��=����mG��t��sQl�0 ��u1�%��;K�Z6�xI���?$NT��P�y�"'��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�KpY9��5�Ě��OY��-��"�h7�~Hw������4tչb� ��o!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���$�2_�u�"�H��RҊ�nۯn����T��g�$2�b�����8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i32e�6��ѝ�9��&n��������QK����ឤt