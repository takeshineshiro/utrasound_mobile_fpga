// megafunction wizard: %ALTLVDS%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altlvds_rx 

// ============================================================
// File Name: LVDS_AD.v
// Megafunction Name(s):
// 			altlvds_rx
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.0 Build 132 02/25/2009 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module LVDS_AD (
	rx_in,
	rx_inclock,
	rx_locked,
	rx_out,
	rx_outclock);

	input	[7:0]  rx_in;
	input	  rx_inclock;
	output	  rx_locked;
	output	[95:0]  rx_out;
	output	  rx_outclock;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: Clock_Mode NUMERIC "0"
// Retrieval info: PRIVATE: Data_rate STRING "600"
// Retrieval info: PRIVATE: Deser_Factor NUMERIC "12"
// Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
// Retrieval info: PRIVATE: Ext_PLL STRING "OFF"
// Retrieval info: PRIVATE: INCLOCK_PHASE_SHIFT STRING "56.25"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: PRIVATE: Int_Device STRING "Cyclone III"
// Retrieval info: PRIVATE: LVDS_Mode NUMERIC "1"
// Retrieval info: PRIVATE: Le_Serdes STRING "ON"
// Retrieval info: PRIVATE: Num_Channel NUMERIC "8"
// Retrieval info: PRIVATE: PLL_Enable NUMERIC "0"
// Retrieval info: PRIVATE: PLL_Freq STRING "50.00"
// Retrieval info: PRIVATE: PLL_Period STRING "20.000"
// Retrieval info: PRIVATE: Reg_InOut NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: Use_Clock_Resc STRING "AUTO"
// Retrieval info: PRIVATE: Use_Common_Rx_Tx_Plls NUMERIC "0"
// Retrieval info: PRIVATE: Use_Data_Align NUMERIC "0"
// Retrieval info: PRIVATE: Use_Ext_Data_Align NUMERIC "0"
// Retrieval info: PRIVATE: Use_Lock NUMERIC "1"
// Retrieval info: PRIVATE: Use_Pll_Areset NUMERIC "0"
// Retrieval info: CONSTANT: COMMON_RX_TX_PLL STRING "OFF"
// Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "12"
// Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "ON"
// Retrieval info: CONSTANT: INCLOCK_DATA_ALIGNMENT STRING "UNUSED"
// Retrieval info: CONSTANT: INCLOCK_PERIOD NUMERIC "20000"
// Retrieval info: CONSTANT: INCLOCK_PHASE_SHIFT NUMERIC "521"
// Retrieval info: CONSTANT: INPUT_DATA_RATE NUMERIC "600"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_rx"
// Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "8"
// Retrieval info: CONSTANT: PLL_SELF_RESET_ON_LOSS_LOCK STRING "ON"
// Retrieval info: CONSTANT: PORT_RX_CHANNEL_DATA_ALIGN STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: PORT_RX_DATA_ALIGN STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: REGISTERED_DATA_ALIGN_INPUT STRING "OFF"
// Retrieval info: CONSTANT: REGISTERED_OUTPUT STRING "ON"
// Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "OFF"
// Retrieval info: USED_PORT: rx_in 0 0 8 0 INPUT NODEFVAL rx_in[7..0]
// Retrieval info: USED_PORT: rx_inclock 0 0 0 0 INPUT_CLK_EXT GND rx_inclock
// Retrieval info: USED_PORT: rx_locked 0 0 0 0 OUTPUT NODEFVAL rx_locked
// Retrieval info: USED_PORT: rx_out 0 0 96 0 OUTPUT NODEFVAL rx_out[95..0]
// Retrieval info: USED_PORT: rx_outclock 0 0 0 0 OUTPUT NODEFVAL rx_outclock
// Retrieval info: CONNECT: @rx_in 0 0 8 0 rx_in 0 0 8 0
// Retrieval info: CONNECT: rx_out 0 0 96 0 @rx_out 0 0 96 0
// Retrieval info: CONNECT: @rx_inclock 0 0 0 0 rx_inclock 0 0 0 0
// Retrieval info: CONNECT: rx_locked 0 0 0 0 @rx_locked 0 0 0 0
// Retrieval info: CONNECT: rx_outclock 0 0 0 0 @rx_outclock 0 0 0 0
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD.ppf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD.inc TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD.cmp TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL LVDS_AD_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
// Retrieval info: CBX_MODULE_PREFIX: ON
