��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�>���U�_�4�0S�����x$.:&R�nU���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍C95^T��6\Xa��7��Į�N��=i�@x_\q��oGo�Z�������/�)��ɖ`ۺ����N<��;��� B]�pE���	x]̃Dj#^Da����M��@D'g��r�� �u�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|����w'��1�:�Ω�>���U�_�4�0S�����x$.:&R�nU���T�����\�4�sW c`k���(�Y���mM+­�\��S�Q�L�����Y�b�Cj�,\ަ�It��vȯq�
� �AH���g���	�'�Wا[b��(�s�J�=�ʝF@�4%���IR.ux'V�vЊ�[-d�x�����q�M�40�W�wƼ�{�4��W��#0��<JTT*��@n���SۣFߞ��G�٘�`�Ocᑕ:�,��JCq��jr#�9l$!kdq��]x��	�VE��t����G�٘�(�����3Y&{ �ŠB�N�M2rӪ���!�Aͧ�	&�~��FjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Q���Ӿ���	���q��q�©�����<�������~s���^��y�g�M)ԉ���S��(�B4�rs�F�r�f�t�B�wj$g�a�\����Ŵ�(??a,����\{F˯�+)��ʺ�;[�ʆ�In��t��Q�]���h�S{�5��lW0��E����F}�=Ll�����,۽���}i�@�5�}�]���"�,�>E��4];ˍH�7��_��To^�|\5muXSr���K�d�eM�bmx�]�V���)</����k�*6[h���	;h�)�[���6зq8�Ј)w�<�_N �VL�(\F�c���$/���i� � �	{��$�`V1����Ea��Z鎬�������(���P����ˮ��lC��U�T�\ ���(�
@��^��1�<��<��z��}�0z�cUL�n����4���á�~O�"j���b7���Øfq�\E��0�ŭ�����]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e�,���6+��A�y�0� 7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7���Øf4%6� �77Ê7�E�4'���Xw�f�VHF��>BH<M�z�]�!����M[��Ǣ����K? T�ҋX����*�QN����q�1Ig�I�?g�f��Qө}�8o�C���7I�����
~�d�9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8��������?9�M�Ч��Dua�\����G7��èV!�����+�yƔ��u����L��>���	��z���AZ���$1&O�.�g3Z�j5�{�CL�x��m_�/��!N\PPE�H�b"�uQ��z/�B{�o
�s��$�Z;��|B[g�� ���S�@�
37�˱�5PM�^-q�x�l��1:�N�*�xSƏw0���D ML:�,�Xʚ@h!�`�(i3!�`�(i3fC��T����ܼY��j3��� Q�N��*lOO_Nc����L�{!�`�(i3,��O^�{	��O� m5Y��j3��� Q�N��*lOO_N�B�r��!�`�(i3,��O^�{	��O� m5Y��j3��� Q�N��*�������)�ak�m6!�`�(i3,��O^�{	��O� m5Y��j3��� Q�N��*�������,�Xʚ@h!�`�(i3,��O^�{	��O� m5��!=.�
kZ)� [��v���Q:�g�a2�-�!�`�(i3�5�9�(��Vh��W��'�u�uX]�Rn\�_�B�r��!�`�(i3!�`�(i3fC��T����ܼ�r����`�4,�pI�!�`�(i3!�`�(i3!�`�(i3�^,�E��HS����ݚ�Н����Y�l,r\����!�`�(i3!�`�(i3x&_FA"���@�ԗӯ��es��O!�`�(i3���gRI/,�Xʚ@h!�`�(i3!�`�(i3��q�Z�n&Y��!둿,��L�������$e����C�9Jn�+!�`�(i3!�`�(i3���׻�t�"hzf�?ǉ�=��4tBu6�]���~!�`�(i3!�`�(i3�X;p`�C��[���ԗ��6%�a���!s�;�����,�Xʚ@h!�`�(i3�&8�,��i��F�ef�?ǉ�=��Wʁ�w�*�fBg�!�`�(i3!�`�(i3�X;p`�FJ���f�?ǉ�=�T55�\H{�U0X��~&����}Y{!�`�(i3�X;p`����ݚ�Н���>\�${lZlX�l��)��40� \��M��ǂ<���HA)��j)yc�n�.�_�t�f�?ǉ�=h�q��d[dͤ���!�`�(i3!�`�(i3�X;p`�;-;*�7��3z%�u�܆7p�J��PW�o#�_T��!�`�(i3!�`�(i3!�`�(i3�^��9R�^Ƒ��f�?ǉ�=��<H��c����L�{!�`�(i3!�`�(i3�X;p`�ct�:��RE3z%�u�܆7p�J��PW}ݡÝ���!�`�(i3!�`�(i3!�`�(i3�)ύ^��R�^Ƒ��f�?ǉ�=��<H��(����O�c����L�{!�`�(i3�X;p`�����L�ҀL���Gk��,�:�N�*�xY��j3���������g�Hn7�(���6����%�3��{}�́��!�`�(i3�-���k\�H��bf�?ǉ�=J�a3mPy��ۊ���<+:0�!�`�(i3�v1a{J��w��!+��^���X�2��}��g��9|P7�_M��f�?ǉ�=����Gx�6_s/ֺk805;<�!�d�<�.�g3Z�j5�{���������ڝr�F`�n��C��ip