��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��U��}��x�� �� ������[���a�8%`��4�s�6�XAoeu��a@����þ�V��1�Wqlw��9�K���m��+o���sp%��X�����b1Ø^���#K���lӧIA�a�V��R�bC o����܊J�j�K�J�'�دv)h�V~�$v�p��"}�vo7k2a��pP.S��*����طǪh��p��U>?���>�`\��Yi���u����l�|���j@��"�O��$� ���xI+r�� 0�D�A�f�mXׂ�(ѳsv�`�S��Y�ix�P�Ra����+��a̞w���{ֱ@�W�8d4؇��2O��'HY-�z����s�1�WNcz7\F���r��RL�a))�kc�߇N	:.���n��{�'��?ɮ��N�7C��Hq-/��@�]\���<��9�`J�=�OLl??�L��y�����c��(r���U�N���AZ��/��aG�k�8���҆�|n��]W Z;��T����G��F��=��J�Й�m����ǥ�P+<�F�z'�_��z�Ӧ�'�b+aQ�wT�	$~j�u?a'���]����Ϭ	N*�b��n.�G�@���y{��O2��@����ا�k�8���҆�|n����wH�L�ƚ��Թ�'�X�׼J�Й�m��/K5r��!����%�������Q���K�u��\�4�sVE34�@d�)����c���w�]� ܩ�*�o?�M��;]�NT[�=� ����i�D���_i��Z��71��%�}Ř&�� �W�#!��Y�:pRр��>�B�m�!=�y����h�}�)���32�d�87��{H������o?�M��;]�`�}��_����Qr�O��C��0���/���k���_0��*�Ε�u���;��.~�Gj'��w9����`e�TS�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����2�C�b��}Y���%�5�1�:�Ω�`<4}��)�Y¹w�yB-j&?��2�C�b��}�{b�2"���Bpш�#w��q�©���B���������'Sea�8���`<4}��(����5�2���[@%����nEAJ_�'��P9��6�g�m��+5z�P�_XV�>!�/�7��u���nEAJ_�'��P9��'p�@�I�?g�f�,�� zr����$l-�㰻��1}Kط��4q�����]V�H7'�R�^Ƒ���E����F�'n�^0o�\<cj�Ur^�R@Κ�2'�̗������\�ݠ�3zL͊�q��UG�s���AE�HÇG�ݪ���[7�d|���XP��Ȩ�wl��h돮h;e��w���U��7�ܥ��2��&������4��5c'�0[����	��N�Ae�#ͷ:��6�J��j��\w��0]Y��
�iC��|g�Y�'���Xw�E�i�m}6*�3���f��]���>����Cη���YL��[�T:nvS�)37J*u>����C��pMݦ�l��-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0(����!
%Z鎬�������(���+�0+�]4��ݪ���CyW�f�t<|����faՊJ�e:[e��mea�8����U��}�o���#ɀ�Om�����67�a��c���}��D���(��z�j�)�q��1�:�Ω��x[,�Ns��{0��d#�R$��O��&�k��T:���V��9���Y��_E��V�no#��٠R�^Ƒ����"X��[��Q[R�7����n9�jsrCm�kO�=�ͦ�ڛ��4W�U����z~��6��	���`y����@����gG�[bGf�ޡ.pz�L�Y�{'%s���'����no#��٠R�^Ƒ����"X��[��&b2��sv��q͆c�!{p85��c���鿋�E~���W�6?��V���>?Mno#��٠R�^Ƒ��e>۵��>3R�d�ܦ)ݝOv%e�Vi���'�)�Բc��j*���F��
�D"�i:�gR���X��O���r����!�`�(i3����}��T��{���ʻ`�φ��<�6�@a� ���N����o�|�B��o��7�dPi��Y��bs��2[�a��o���Pi�#��R2W���R0s��>H�,b�z'hۉ)8D;�:㰻�߆�p�hؽ!�M��9�a>*<UB3 �~k�%�����Fodً���Fz�e<�Ia��la��o���Pi�#��Rq�\E��0谯n%�Z�'���Xw�j�7��+�uB;y��.U(�HN��R��#�mo�����Ě���R�`�)n�S߸��S�Ȍ`�*Ft���r%k$J&+��T�����D3���������M�ϸ��#|S������3[�u8�U��֜��3!�`�(i38!�w� x?����,��L��$Q
ˋ!E\1�1�ҕ-����M���R��ӟ-����6%�a��'abW�5�}�]����x�8�D"��a��'�-�H#�"8��jo���po�h0�h�#"
s���
|�1�0j�$��:�e�h�Ϧ^c!�6 �ef��BA�IH���O,8��=����t�F�,�U6�Q�L��֭�h��O5�tx\s�l.�	�C���ɕ�eY�����w6YmC,igu[�л���7M+э4��Y�{'%sd���8tjsrCm�kB7Ԅ��p�n���d�)bU�k/9$0fp�m����&k@C�Ɨ0z�cULb���H��U�H���3Ah	)ޟ�I.��^�