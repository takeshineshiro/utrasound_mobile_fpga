��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�L'jf-�6U�P�H�q}��������]��;�Iώx�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R����h�K�5���� ��1�:�Ω�=A���>�L'jf-�6U�P�H�q}��������]��;�I�����)O��Ξ4�"�\�� ���K�O�{����ۤ�9is)V��㝒c\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<���-ZW�k%u�e<��⪘����t�켻�S���c,� � U�rN�3��m-�@xI+r�� 0�D�A�f�mX��VNF��SK��1�����o�T�Y��6�C�-B��<���2O��'HY-��Yk"1/р�{:��'��팣+����F�N~Y*z�w4G� ���������	x]�V�����v����,B���_ġ��M�S�O1��*F=ॵ�h��!`Þ3�����c���.�6X�,4�?n5���AQ� ;-]6�*20��K�X��=o����"���	x]̍�9��H��@N?�qt�-U��S���D	��e#�'���'�A�n���Bu����\�4�sƐ�hd	���Z�<uoѼ�=nq���i}3�L����­��+X�0�w�Gu������	��wˏ����J�2j���_��J��RL�a)'r�Ӟh� �������JܠR)1���;$�� ֹY���8hjY탌�S[W���9��1WA"SӠ�|&�q�!h���噞� x�����Kr4��n�:��e]މ�;���J�	�هU7S�>
��W�Qx�ـ� {�����G��D��;B&�� �=�?��"�Tp!!v*!��1�����f��{0��d# c��(�U����	x]�fX�eϝ(�&Vi���ܩ[߹f>N�u8t������kk��������yȝ�No��>���:E[Kڱ�cTm�Q�����<D���Yl�2���[db���"�p�����J����R�"+���Ŝ�g���
� �AH�W���,v����,B�_�>��\�A�D�S�O1����l�n�Zl���H��6֛Q��RP���敿���|q.;�aE$ /j��sZ19(�?Z��pV�����U-�P�?��ԭ� � �n^�*���j�Ƿ�:h�(n c��(�U����	x]�<���e���٬���f��S���D	����,R�/�G�m!7�X��@$W�ػ��Y�׍�C�	9�/{�ڌ%|w�u�]bu̎}�Zq��Ь��dy�D��3	�53�'6��
�U��p騥m�!=�y����h�}�N�5�%���3�3� ֪-H��U�)��NT[�����=��A|����n���g��k�8���҆�|n����0ӵ�q�TGWXR�� �*xf�+���B�x�
�b+S�������\�4�s��{��]Qǯ������(2�SnFUR�.�;�~�MUs �9�N��U*��$1Xf_q[o��>�`u^9�렕4��S��$[��������\�4�s|��Z�w�N	:.���nњ�@I�y���޷����7C��Hc)𡔚I<Y�@�Nq"Jc�l�!H���uS �����g�Y!#v��v�0gSx̏7�ɍb�e��}vh�xC��6֯�x9���z�{AN��L��xScKE#���,��n��zWi@�!����,x�}vh�xC�}��C�p �Q8�m���8��!�3".t�|6
~����0_�r�O��C��0������m�Q 0��]�������n�u���;���A��j`��'�����`U+n%K)��k��Ǣ���N�y�Yc���;��sD���L��+�Uz�QLQM��S�O?�4�ʗ
� �AH��1����̷f�R{7�2�,`)�
��5i�ĞX7�F@�4%��"�-;��h\kY��%4]��4l/4����"����U��y�Zk�Ž��=v  [f�8H��0�0�G��?�d���&�3�S��3Ze�P4��
� �AH�P����w'm'���h$4����3�^�8A}�؝F@�4%�}����b�+gobQ�e��R�-9�m�!=�y����h�}�~߈#����xy�V�YP��0)i�p&�K��~�MUs �_ܽ�Xr����7�C�p�e$D������qθ��=D-0m ��Q����=��u7��
�+�0����rm��?�X�'2)8�6޽6�H3����1��OV}�L-e �Q�����qθ	J�7-"8��G�(��k�8���҆�|n���eξ���k�o*1��b�T׿s�esP��F@�4%��2@76]\�B( (c��G��Dv�EO�{���4[G��P.!܃��L~΄gO�3T&�r�?^0�f�W<N��6I�"�B�Z�Ӛ%K��SQ�B1�	Bc	{���C<G�m�!=�y����h�}�)���32p�D2]'�h����%/�o?�M��;]��,��K!�n@�{IT̽ae���m�!=�y����h�}T��nJ8�TT	q��$a4������LzX�AX�~�MUs �ˠ{�t!�.�r�c^�e���zǒBs�&���b
� �AH�T�t��3��e��ME
^����c�:���0�F@�4%�u�L�r��3�jT!�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3����M�	g�y�+��T��C�NJ���1�:�Ω�A��>s>;����M���^uq�.�b���q���1�:�Ω�S�T�;Ϗk[�^��_E$ô&y����c���o�����0�ea�8���	�~�����F��mF�!؂������uq9����ea�;y� ����t����M����3��~ �Q�^�y�zL͊�q��UG�s�����M����V�܄WD��|�����u*K6HT�����N�t�&_���9�!�`�(i3l0��F��j�q	k���Aj޽���Ǜ�����������i�l0��F��jT�����N�~ `�T�v��1��B�wj$g%Ah�%4
>��XP��Ȩ�wl��h�d�uY�؃�]n�� ���3�ҺIÙ=�H��ˡ�VkLs��dJR�^Ƒ���Q�^�y�zL͊�q��Yy�u'�7�;�r��0I� X�1��E����F���8�TP�}{�Z
M{2jR�j���m l�o�����зq8�Ј)w�<�_N �VL�(\��'&S�39؍��R��j�.(Wx*��|��pe���b������5	���]���>����C�h�'f R!�`�(i3��|g�Y�'���Xw�E�i�m}6�B�r���E����F��j��\w��0]EOJ�uxm�3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_��ct�:��RE��W��_�ړ8���/��^����r��H�+k&v�Iz��j���'b�t	�U���C��O]r�<Uee�,�Aٺ�H�NI�:7�N�5�%]���a(􆿳����)T������ݤ�v�ϭl�\ѵ�Th�fܯ�ko��o�����}�ꢤ�OgZ)[���F�����E��@IE�U����S8�����NlU����z~��6��	�\�HP@�a���н�!	ozqP�"B��$I��w��,�������ݹ�0�������Dɵ�p�AJ�e�$��\�*P���8��';�¬pX��g��U-�eaԗ5��C�6�ǌ�lA�1�:�Ω�=A���>�L'jf-�6U�P�H�q}�������Wa�b����y�E�nwE��S��}|��XH�����,>$+W��� j�(����5���I�zI.�R7�$��p�S$�&�R$��(��]�/(f�|��*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e���b P�|h{�T��`�)�	�%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��Vx�%L��W��_�ړ8���/��%���aX[�=�5x�� �i�#n����Ր�z*���Be�2l��4��a��se�ξ������ei4����/��)}���/��r��H��p8�(�E{p7�j�pܔp�l
d�R�.��On��M��ҹf�f3'�YK4U)	��$��Xo��yذ��t�H�MPq6.��W0i��^%b!&��曯����P:�UT�P>&�&i��w��9+�7ޚY㮭6��.��LLn��S�W�כJϾ�i���8��'������Ů���zO�fIZ����b���=:Ln��S�W�
����uK�����.��4�F1��������ň�� k�|6�8��^5(9�։-�.l?e�>����c_����+�˂߮<ur�<Uee�,�Aٺ�Hۄ�2HG�T�gs �\1�Z���=�"j���b7���Øf}�
�?�?KYC'v���NE!/��Vh���*ܑe�W����n�4�{lGD�V�B��иܖ��A�.u�r���,DTc�~y��i3���w�@V�c�x���H@H�֦g�㎏qló��@d���/��=��K�R�hE!3�͸@����gG�r�I��!�`�(i34K�)s"e�>�������e���"}�`�W��f�(d0iV�6IWJE�\��[�B#���1���Q��ǺΕ������5|��>�N�B��3�>�>���%���e'6���;8=�g��U-�e���b P5b11��m$��O�&��;�L���9��Xv7�j�<���dW�ML�f���m���V��_�Ps�S��u���2ا@�����ۥ0J�G|�F7�_���|�Ya�ь�+����eǎd .8Cm?��>�&n��{Xm��B�.辪��|����OxtX+�Y�S��?��L	�<���BSz�R嗞Y�{D{��?��L�de���"�m���r°������R�wX����K�Q_'&�d�'f�lR��~�ό� �������g�[��w��5�e`��9x�P�$tw��z䮃\w��0]b!��u�����9�H��@�Y�:/��N��I7��-5��6��	���`y���pzl��a��ҕn�s�� �ߎG�a�x��{�6�e���ӯIJ ��`y����@����gG������G t"���ȵ�ixUS�o���ia���lC��U�T�\ ��i3�|)sՀ�/V������?��;!�uSP n��"(ߔ���?��5�%]���a(􆿳���Qs����� Ei�lmZM������)��Q]� _�rs�i��<�M�AϦ6��.��L�=��gr(��������B�D�F Ho}2b<�TC��G���-o���Y�{'%s�O��W���"�m���r�{q-Tjo�R�wX����K�Q��x���!����a64Z鎬�������(�����9x��p��;mQ��8���/��9/�*0�`R����}tm+�͹)�"�vҕL5ӥ����S�ۗ�	ͰZ���0%�!�7ӎ�؊�"�Dz�Q��y��èV*�n�'��9G�#,��gR� �ұ7���?�!� ��X�J�RgR� �ұ7���?�!��Y���B�?�9�e�Dcb��܏� �� +@���,@��y&�楰�m l�o Z,l��lH�r�hr�W�j#�{D�A������G%Ǐ��� gWVbT+zv�؊)�x��d���!i�RɆ��_줧F�5(��j���rz+��bc�n7�}�!��g_��T�d gWVbT+踫g(�r� k�|6�8�Eo(d�J��:����5s���Z�����t�T��?E-h��$^(?��"��K��O.C��ݚ�Н����"sS<�0�zG�������&G!�`�(i3EOJ�uxm�3���w�@V�  ����'K7͍��|��W&":�ݚ�Н�ЈH����@�/�M�k��G<Y�dN�<@Iv��nt=:��:5A��p���aR�!�`�(i3�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}�����l��=�O�-v�*_�mS8<�n�ݚ�Н��wӨj]h��_--���g|�m�ߕ�v{��lw	�����4�:5A��p!�`�(i3�u��g��L���ʗ�%�A�i�A�r��H�!�w(�y?!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �W?�;�끣�os�鮊R�<�t@�.�g3ZY�T5��܈��zNc5�V��	��y��=-f`Rg.�YP�׀A���`����oȺf��m<�E��?�d���&�t�{#	�x��_--���g���R�?KYC'v�����p�*��nސ��3���w�@V^�h۾�(z�k��E�2}�	76�&�;��|Bת"tg �+aT��3G?�d���&�ϪE�smy��]=c�����<�g�daBb�KM������p�a~�'�� |X��|̃?�9�e�D�a~�'�� 7��
�+�0$��b��{��2������<�b�)��:��?�d���&�C#/<���q�<��>���-vR���B��G���S,��!^·ʌ�C@�/�M�=t�z 7�J�[�?:ͪ�'����,�ǰ�L}��t�gb�"�?��A�rD����}��\CB��u�Y�KG�	�v�3� k�|6�8��:�EB�Z5�O�%E#P��k����  ����'�W�6?���_--���g|�m�ߕ�><���@��`.��53���w�@V���<��I$��6�F����������o��_�Rv�䩲$���dS@Ɵ�o8����z�(����<m5��IM�Ex�>�+X�M?��y�!�`�(i3�y�, >����صW�my$�N��o�/���;�� л��Ro�G/]%�z�-uͺ�s�η3G��Hb+�����;y��v��\���
^�ݚ�Н���fCI��8��GM2�]�<�k��u���H�����0�و�@Q�kj� �v�қp �F��ݮsȸ�"rR-��ټs�  ����'Z鎬�������(���kO��u��<��>��h�EtC�<����J�F���i���ϴ�����?�618�V�
�>(Z*��b!�`�(i3�Y�m�k?j���Fz�8��;Yv^�-w2M#-5�]�!��	Ǹ�y85��X��I�ՠ��t����>3���w�@V-���,W��AԢ�a\��MԵ�x3���ʗ�%oc�����k��u��fĉ>99��A0ok�²��y��lDX�t�VC��c�{I��L�1p/-�������?�/5��"}�a�x�mj�B��Vh�EtC�<���v�9�ʝ�\ Nh�;�P�t�5�� л��5ߧE4�흔\ Nh$�)�vx��������;_��8W�w��fD2�es~�@IL<�	��V�/�z�r8��	J���6Oк(cJ��\m�Q�  b�ۋj�[ʙ{�x�۶�kv�ѓo˄.�E�t&;��.u0B�r��u�Y�KG�	�v�3��<ͯ�G��R'),��`�a"��-K8?�d���&���n4s1�+��uK[F"O���%��ɶCmsW�C��`6���ҹ"��s��?%ww��Q��ǺΕ�=Y��~K?�d���&��ݚ�Н��9�|���l8�48�{.S�����g��+˘\5���jmY�wΦs� ��6��.��L�la�F�wF�,'�*;���#�b��{�.�t#6��.��Lj�)6)-
FkH���8ч����B;�T��Q׭n�L���/=9��9����C.�L:,�s L�Zl�W��{��]�L���/=9��<��&C.�L:,��i���A��;b�-�2�V��	��ypw�|F���}Dq�f�R(��N���v��T/q3b�5*s6=��GZ>.�0'j�j�Jy?�d���&��ݚ�Н��9�|���l8�48�{.S�����g��+˘\5���jmY�wΦs� ��6��.��L�la�F�wF�,'�*;���#�b��{�.�t#6��.��Lj�)6)-
FkH���8ч����B;�T��Q׭n�L���/=9��9����C.�L:,�s L�Zl�W��{��]�L���/=9]�5LdW�Q���=)8�+���LQ��:5A��pw�R���y��[�ڰ�����"��L��:v(ȉ��G�
Rv���'\://��=��K�R��K<_8 _��s�֙7�}�!��!q��V���'�Pp��XO)�Q>�W��*(��3H��ieL���1��#��{�6�e
��>�i�g��+˘\5���jmY����A�I�{�6�em�;���Zt%��m&<XdYʼل��OY'�E�g�������(ӈ���m�r����I��)���W�w��fDC����^\���b����	�.8����-��1�&l����$�<�F�q;��|B���r��������o�a�NO�*b*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���r!|�α+SƏw0��N�ijR2t�N�/�ڂ�nF���<�W�.�P�	��
�Q�}�.�g3ZB�ek�5W��x[Gň�����f��2Lt���U��)���Y;e�iKI/B޾PԐ#��go`(&�L�xjzӝ���I(͂��-����Zt%��m&<o~葸ֿ2Ĝ�sdN�<@Iv��nt=:����q��{d~~!"s�3�)��b_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:���T8��Ʈ+ˀa��z��2�,�s�Yls��8��GM��-����!�`�(i3��8���L��Z�|�� �X?�V8ч����۝�n����Y�VQ��$��v̢����9�|���l8�48�{.1�m+�D8fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx�)���+��%�q(�_��G=X����>1Y�V��	��yv�ʯʗYo��g����~�'��BP+>B@H/b͠�Ԏl�Б�����ph�)':�f-�Б�����ph�)�w|�0)��]��.e�����م���R7�j�2>n�IՏ��J��:����2Zwz����1 ����C�#�,�IX0F�MV�ҁGG`5:��"�9ŭ,iI9�o«IX0F�M���`3�JV}��� �I!�`�(i3���{���#�0�zG�������&G!�`�(i3�iڈ(��֟�z��n�*�&�v��K7͍��|��W&":�ݚ�Н��B�.�4Ӭ�P8��PS~B;�T�dN�<@Iv��nt=:��:5A��p�I��Yq0�ʂ�j�Ï��	�l�lM�3 H�RtV�^;�E����=�O�-v�*_�mS8<�n�ݚ�Н��� л�������b�� �_&l����ۙ�Wl��pH�RtV�^!�`�(i3�ٻY84����<	s/S�����g��+˘\5���jmY�wΦs� ��6��.��L�la�F�wF�,'�*;���#�b��{�.�t#6��.��Lj�)6)-
!�`�(i3Z��}	���C�ݥc&�̢���>�W��*(��3H��ieLb)�5�o�' ���@�0�0c��L>�W��*(��3H��ieL���]Cr$' ���@�$� %7�!�`�(i3��\ NhA� ��_����{У��иܖ����Sp��;�{��!�`�(i3<�6�Q=��hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]vK��L�'`N߼�K�iN�� ��t΀�+I@L>���@]��}Dq�f�!�`�(i3�ٻY84����<	s/.�Ss�g��+˘\5���jmY�VS���g�n�{�6�em�;���!�`�(i3�^{T~H��������>vD���&l����$�<�F�q��-����!�`�(i3����j��`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3<�6�Q=��hY-N�g3�)��b_X�XV�b�z'hۉ)��d�7�q�!�`�(i3�^{T~H���r����!�`�(i3�ٻY84����<	s/S�����g��+˘\5���jmY�wΦs� ��6��.��Lj�)6)-
!�`�(i3Z��}	���C�ݥc&�̢����{_8�Y��=�}�Vݨ��}Dq�f�<�6�Q=���F��O��ݚ�Н�0��l!���O�D mWN<�6�Q=���F��O�ȓM�Me���]� )�+�~�8�r\���1 ��b�i3�0��l!���6j�"Hs?Ճ�1a.�&�"M��N?�&�{C9	��9 �l]'\gWg��	�Z�kfc��2���8���+�^U�	Y���xjzӝ���I(͂��-����Zt%��m&<����Tif���GK7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3e<�Ia��la��o���H�RtV�^FkH���t��@����Ŋ5�m�o~葸ֿ�|gԁ~~!"s�3�)���:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6������}��;.��<񪏧�Y<��w:��<���eʣ͜��O��a��nX�������o<|O�Ӈ�t��<ͯ�G��R'),��`ޢrA BG֞�"'�Z��
������o�C��f��26��U��ZW��:�nΏ��Z��L�dGk�>}�����L��Ay46�o8:4�I���c�90�Ǘa��xO.C��WHe�Q\���F�`yx�>�+X�M?��y�!�`�(i3_'&�d�'f7��W��~�>� {�}���my$�N��o�/���;�Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#;�jmT�#�,l����M?��y�!�`�(i3�#~.��,!,�:�� ���?R ���8����]�����q�w���팣+��!�w(�y?fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��.��vذYC�8����g����<�c�����M�~���!��w;��P�{���zG�b@�d�tO�+�Jam���)�/��� ����H�ʱˡaf)��S7���8�K�����.��4�F1���l혡˻|��X:< mjR}���܁���e�[�O����� ����H�ʱˡre_���G;��|Bﻍt����-�����#�Y�Cφ��<�6�@a� ���N���������y��o��7�;�jmT�#bs��2[�a��o���H�RtV�^�#~.��,!,�:�� ���?R �K7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3e<�Ia��la��o���H�RtV�^FkH����T����!�숫J��M-03�gM�¨ɢ�=��g*�ݪ���c�0��:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6������}���팣+���������V��	��y���"��lH��H"��Th�76AyW�Dw��V<�:]���7�nξ������QNx��f%%eTe��`����e����u��.tƁ��b�������J����;�f62,��}�Hy�'9��ł���J9ߝƊ�}=�s)��!�VMJ�KC�}�R�۷���z��U������>���c�m� ����\�Q��4b&��K����8��ۉoo9��#U���Ʊ�_�eD�I�6Sa쎑Gc~�;�b���=:�Xb`_�yK�|q��=H��6���,���eFz� �l+�8�#��'J()������TV�������j;�㡙�6.HY'Q�w��������z=q����\����C9C�!�.g�e58=#`���g�W�2AK�l=�"v�(=?�w-��U��)���Y;e�iKI/B޾PԐ#��go`iI9�o��|#HK��A(�c���_G��Hb� h�ҩ�!q��V���팣+����ß�m���nF���<�W�.�P��c3��ɮ���Ł����p�my$�N��o�/���;�Ra])n#�璓�c�������t �[l;[�G���KlG%��`��ǚ��ظ
��@�U#;�jmT�#�,l����M?��y�!�`�(i3�#~.��,��tE�ӻ���+.S=��!���c�A�L'%=}�^�m溼팣+��,@[ܬ�c���k��$(�%�8��@�A���Y�VQ��IچG{��]�!��	Ǹ�y85��t���]gM�¨ɢ��9x��p�5��/��8���/��:5A��p$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6������}���팣+��#���@���]��.�Z�eր�����,JjH��1�:�Ω�P�p^��J���t��������Mt�iZ]XF�hx��G����Tkd�_Ji�];���Q��\@
�Q �H����]g,H��vє�&���X����?����O,87WA��s�E���g^{ʓ��(%��A��)�^�\�E	v��o�1Ʌ�Mi5�'�@b��Oa�@��I�Y�K%-H�V�;���)"������w6YmC,iguGظ0����t�%�Z?�MZ�ʛ�z���dЕ�ĦsW�0�c��,�#���@��^{ʓ����-�����<ͯ�G��R'),��`�K����F?�a�x���x����A�l$�+9@[�_zβrE��g�Hbc�m� ����\�Q��4b&��K���w�����z���o������,�ǰ�QCT�"��I�N	�7Q�n��;:��_)�:)f�����9x��p��;mQ�MM
��,=�GdC�b�>y�T�.�~�k��D����팣+��A�׭�%*be��0�U+�qbp@��-��~U��j����J�;����<�����;�)R2�bP�=�ƛ������CyW�f�t�}+N_q��(R\֎u��Vv/�y��{pxʟwf5��F�$N!U�t|�Vx�%L��W��_��MM
��,=�GdC�b�>y�T�.�~����`���ƼP��d�k��԰�/"��nH�W�q3��+����/���	0xǎ� 3�kM=/[�)�������sP�������tw��ĕ[뜗��,�ǰ�ƍ��i����E�p�2W���R0?�@�|��Z鎬�������(���R0�����%��Y���#�����.��4�F1���Gb	l�%T�#�S�� n`Ip�\{ف(�7���<��Y�&l������8y�Ɋ����Z���F%�X�ԼQ�}�p�?7P���`$�P.eE������v�h�g��U-�e a⣃_B7�}�!��?KYC'v1��E:z�'�=;v�����Ə*J�X�$��c��GlhŦ�.�g3ZrZ�0m�\�S��u���F%�X��/����7Fk����PqZ�o���ia������v�h�g��U-�e a⣃_B7�}�!���u��g��L1��E:z�'�ĩk(�CQ�r��H�*J�X�$��b���9C�.�g3ZrZ�0m�\�H�z��.�g3ZE��g�Hb麭�H�κ;q�+����Mgw�� 
~�F�,���XF:6/������,���eFz��^�̷ؠJ��:�����0c/��kk��o������"O��_U)�<�&#R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P�G��^��jsrCm�k�:��=#��9f2Pih{Ø�Fɝ�\ NhV��	��y�� �P�qN�/9ݦ�R��X鷴QW�w��fD�W�_����Rr������%�<�$