��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��maC�S�s-\gf�N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��d�Ƽ(��h��mo������f���F*�#C(��$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us��n��/�FI���O8�yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\�v�{K���$uغGgt���Z5�0L��t�켻�S���c,]�i,ev.,u���z�����>O!����Y�f��a�Z��Vv�c
�����R��Y���`z�X���#�ӓ]����?6z`D�EcX1R_t��z����j��Y�uvr[�~[�#�X�O��P?;OK�BB�a��ރ6%h`��~��.d�o����m7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3t��v'gn�]o��in�m��+�Ƽ(��h�R$��Ct�z&��ÃlO ܅dxF���u$J��<
DN�%Ah�%4
>��XP���C�&NJ=رx���9pk�o��jV�{+��]n���b9����$�n������ л�A�.�hQ3'c���������n|���띂ii�4];ˍH����Ү���/^�yQA��c?A���$v^�1�N�Ae�#�k/�z�xEQc��Et��q���U�ЂDa��(;�A)k�e.��xu	�>��l%i�-��9��稕v�ј�"��Z鎬����$oi�~ƴ<�6�Q=j���$5�?� �٠Fd���e�ш�_(x��`��|g�Y�'���Xw�j�7���(}y���CyW�f�tR�wX��q�\E��0bq�Z��T�I��w��,c�A�L'z��0N�7;�¬pX��g��U-�eE������(fx��V$�w�I�?g�fl�NAS*>�m۪Y!V���g�uE�EYZ/�h�@�o��I�?g�fl�NAS*>�m۪Y�%0���iI9�o�L~΄gO�3��|��[��.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc%�����I���%�L&�{�(=2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�R�Q�XL�^u˶);ċ�L��Vy��H��w�1T����NGq���ÌL��j��5�O�%E#P{y����M�V<�'~1>��v�&[�v �R!��(㒖�����o��_�Rv�䩲$���dS@Ɵ�od�G}%����3f����%��-acwIt�~;�jmT�#bs��2[�a��o���zM#��m�!�`�(i3��4h�=Iz~r��V�n��dK�����fF0���2��}��e�g��)$�{_8�Y��=�}�Vݨ��}Dq�f�����g�Z��3��a���!@�f")z.��W����Q�Y�;y��v��\���
^�ݚ�Н�:
��x�{�\��N�Ś�-����!�`�(i3@ E���߼WaU�?2����W��_��	h����QR�^Ƒ�Ӎ��t,���~��;�,
�:qEp�;�P�t�5fĉ>99��A0ok�׹����/m�����c��aT��3G?�d���&��R!��(�J�4�Ur�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�Q�4��c�T`��.�&Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h'7�T�f�S��J��=���8�8e[m��PC-��i0Q�͹�Ɩ,�m�<��+x�V�}�OiI9�o�?�d���&�S�@�2�e��}@��)�TT�"eZ�Њ7."t�o��_�Rv�䩲$���dS@Ɵ�od�G}%����3f����%��-�����|#HK��A(�c���_G��Hb�8�u?��I!�`�(i3�d���a؅q$��.��m�f.���G�?v��� �+��R���wӨj]h�7M	�\�dN�<@Iv��nt=:��:5A��p*qA����6\�4�@�� �-jېI�q������ л��E�BS�+��U�,�P!6���r�����$XR�QܛOcOZail������&G!�`�(i3p�n��v{��lw	�l����;�¬pX��g��U-�e���B�/m�ڨ�hծ���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ą���%��-����aT��3G?�d���&�S�@�2�eɢ?��x��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��{����]��a8&N C^2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����N������s]?%��h�r�Bi�v�V���;AD�
�N����wvA�qS�F_���ٱ'W�w��fDe{n���nM����J6«IX0F�MV�ҁGG�.Mm-;�C>��Ӛ��S�J\7fF��v�V�2�~�xjzӝ���I(͂�'�ɳ��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3@ E����x����E2b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��?u��C@<�6�Q=��ž�Ć�T���7X���c�}��
�t��T&��ۥ`�[�G���K!�`�(i3�k��M���#�a�Ą]v1�_ُ=9���Xi�X�����j�5�%]���ox8����)H�RtV�^�2��}��e�g��)$�]�!��	Ǹ�y85����[��蛫���dU����z~Ao��m0e9�Q����0�&�����ݚ�Н��̢k����a�x�l?ud(�F�Їj��ݪ�򈟄濫�L��� h�ҩ��wӨj]h�7M	�\���!���c�A�L'M�M˫ɒ}�+@2l2VQ+�3yK������v�h�Q����0�&�����ݚ�Н���w�w:�!�`�(i3q�\E��0A��6U�M�Fqɔʍ1�Z���=�"j���b7|#9���!�`�(i3���F��O��ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끶���A��'#b�i,n����,�ǰh`���i���H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����1�~��x��sq=���#'@Nw���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�r1�:�^��1M<���8���8�8e[m��Xd	�/I%L(Ρ����
�N����wvA�qS�F_���ٱ'W�w��fD|/%�- F�z16�5k����o��_�Rv�䩲$���dS@Ɵ�od�G}%����3f殚z�hJ��#t-|������"sS<�0�zG����ZAL�:!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н�p�n��n��>�my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	�����y��lD�7m�T��Ʈ+ˀa��z��2�,�s�Yls�<Ԍj��_�mS8<�n!�`�(i3�k��M���#�a�Ą]v1�_ُ=9���Xi�X�����j�5�%]���ox8����)H�RtV�^�2��}��e�g��)$�]�!��	Ǹ�y85����[��蛫���dU����z~Ao��m0e9�Q����0�&�����ݚ�Н��̢k����a�x�l?ud(�F�Їj��ݪ��eL���3�1tSjv�!�`�(i3p�n��&k@C�Ɨ0z�cULE��K3�jާS��m��X�����j�5�%]���&�gl��1�Z���=��n��I
�:qEp'{w#/ B!�`�(i3@ E���߼WaU��xӺ��-���lC��U�T�\ ���:5A��pfĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx�HP�ƎѥH,
��X.V��	��yƄ����vGЊp�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ������
~[�#�X�~̬̙�m��:[�#l�O�֧2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�^�wo������me�k���e�Í�x���"x����O�r�1�B,X���q�*��a�ur�V��*s�}F'�n`5�fK�3L��'9!�`�(i3�� л�������@bpVXR�CpE��:���~���Q�W�����a�ү�`���;��|B$�g��� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc>-��n[��u٨p<��K�<�c��=��c�c�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~'Y��UY-%f_��m����ϏQ��8'嬘�����v�h���h�99S�r�F��
M�,!hޖ�A$�P������5d�`UNP�{y����i�q,?5q�w��.NG����Yk���'ž1�|�'����z.��W��!�`�(i3��4h�=Iz~r��V�n��dK�����fF0���2��}��D�o�&��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h�'�ɳ����Q�Y�;y��v��\���
^�ݚ�Н�:
��x�{�\��N���'�ɳ�����aR�!�`�(i3�:W]�I-�G��Hb� h�ҩ��wӨj]h�7M	�\���!���c�A�L'0#P�O�Z�d-�~EL%�G�b��6��	㎾��;|�5�%]���U����z~��7��:��}Dq�f��	��x��ݚ�Н�?V��j�c]���I���-%f_��m����ϏQ"j���b7�S
��n@V�� �9��1�Z���=� �o�XÉ��%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}���,�ib�2��~v�VV��	��y�3�&A��S��V1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��B+<鷁�[���?��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��|=���ac$Ѕ����n|�p[Y���"��㥮�{=�
�N���2�t'�0a�����S2�d�٣���$u$Yo�K!�`�(i3����v�E��tS�$bnN���+�^��BY�B�3�&A��S��ƫ���v{��lw	���:�(������v�hz&v��\��v鋮�����U��)���Y;e�iKI/B޾PscX{�X!, ��b�FP&�ʅ���h7s�9���oL$�����//��kOT���+�^n=\f�5>�j%���=r�}&xjzӝ���I(͂�'�ɳ��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g!�`�(i3@ E����x����E2b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��?u��C@<�6�Q=��ž�Ć�T���7X���c�}��
�t��T&��ۥ`�M?��y�!�`�(i3��t#�V�g�Tԝ��}Dq�f�5�����}Y��	}�@���	d=�4E���b=R�^Ƒ��N���kb�r!�`�(i3��B����U��n�n��)@�])�#����9!�w(�y?
�:qEpCt�w#��@�����!�`�(i3)p �K�b~*��s��ʅ���h�'����u��r��!�`�(i3@ E����̷_��yC��S8�����ZK�����aٔ^??2����W��_��	h����QR�^Ƒ�Ӎ��t,��SX�4/���:5A��p�Ra])n#���r�����2��}��e�g��)$��K���f�(}y���CyW�f�t(�%JvP�X_Gf���D�ݪ�򈟥��P];�
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹�{��N�i���?�sh�w�R���yh��7�S+��M��+� ���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ڨ;�	��o�����C��c^�.2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���m=��}q��~�_1�HbvI�a�L�������	��
�J:���⶷x���S�A>�qF>:�����KCw�6� .{7s�9���o`�-9v��!�`�(i3�|����*D�WT}�
�?�uf���I1d�|u:SQ'���XwM��%�p@�X����t+Y�?�\�W�GCٔ�*�*s�}F'�n`5�fK�3L��'9!�`�(i3�� л�������@bpVXR�CpE��:���~���Q�W�1��	!��[�=�5x��/���q0�W9a!@�0z�cUL�BJ��VR�^Ƒ����"X��[�w�����!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3P`��dpfV����1����	CE��'�$�}�pI�&5O���F_���ٱ'W�w��fD��m=��}q���}����l�����G���5�%]�����,H/��� t���}�O��R�^Ƒ�Ӎ��t,���_II����7����8G��5	�ƣ��6�o8:4�I���c�90�Ǘa��xB��򨙉����D�Mg�{HZ鎬����Ĺ#{��ݾ�9J�ciI9�o«IX0F�M��m=��}q��!����H����Qw�c4~Nr_�mS8<�n!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+{k�h�+P(�	m#�x����E2b�z'hۉ)��d�7�qć�p^͍���5�ź�q9+t�}�;b�-�2�k+Q�h'�Ȝx�5W ��̫(�8�u?��IlG%��`��ǚ��ظ
��@�U#;�jmT�#��"����G��Hb� h�ҩ�_��F���������;G��
̭�!�`�(i3�ʅ���h�����C��ݚ�Н���=�gw�⽒��5���=\�gL���l�5�%]������	�|��!�`�(i3V/loo4#����F	j��25����K���f�@�VҒm͉��%>�rG40�RS���$
�)!�`�(i3�3	{����I�^$D���5�1q3�;�*5��P���<��~�
]^��Y:�����������y�Qn&�ð��T�ݚ�Н�?V��j�c�/���q�pg��B|��rs�i��]S���D�'�)�Բc�<πV��;�¬pX��g��U-�e�(}y��YmҐ�̓=�^݊1�m+�D8
�:qEp'{w#/ B!�`�(i3O�L"|�#�h\@�-%f_��m����ϏQ"j���b7�S
��n@V�� �9��1�Z���=� �o�XÉ��%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}���,�ib�2�y�v��.Sb_�뉺�p�n��v{��lw	��a{7?TQ�g���F��帵6C
�ɑ��U�]-��	z�{�eM���)��=��/�Yr<���5�%]���a(􆿳��jV�{+�K�$ޘ~��~���v�R��Ǭ�e	0��c$� �顆� Kl7�� $n�@ E����[� �_�+\н�+�k�@��?��9)���9a��=��s�_1�⶷x��݆�TlL�_`\G��.��l�N*Cdr�������G1T3��B��Z�>)��چ�^�RtWH`��PrmX������,s�jK`��D�;��T~q�������@��tW˹H��Yw�7DpA�tA����rd@��W���i���L9H��wJ&��WB�*����^�J�z��R�>�c�>Z���X{)��K�!�fh����G �U�'1�Wd��&��.�g3Z�7�4��~},��� �M߯�Px�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���܁�c�^{�$��-y$��|��1���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Q�6#j����$G1�O���8�8e[m��! ���ÙK��<��?�d���&��@����gGJ�y�b[s>Z鎬����$oi�~ƴ!�`�(i3R炾z���9H���qķB�W�����_^Ys�
��U�|�R�w@n	��d�٣���$u$Yo�K!�`�(i3��$W��?k�g���&�<*|k5*+��A��:�0������.U*j�=���F_���ٱ'W�w��fD�c�E�dE�e��	��!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �:�S}����ق���Բ����-��6�+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc8���8��v{��lw	���:�(�V�� �9��1�Z���=�-+��B�G1X`��5��K���f�(}y��YmҐ��*V�M��nDN-Y&yo�q�%g�῰ ��E��φ��<�6�@a� ���N����ݚ�Н� ��b�FP&�ʅ���h7s�9���oL$�����//��kOT���+�^n=\f�5>�F��)�m���.�]��;�jmT�#bs��2[�a��o���zM#��m�!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}�q�\E��0Ww3i�|ł�nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h�'�ɳ����Q�Y�;y��v��\���
^�ݚ�Н�:
��x�{�\��N�Ś�-����!�`�(i3�(MXdvm�QA�Q* !�`�(i37�%M��أͽgF"?�(}y��YmҐ��'�V�k5j[��(��!�`�(i3��t#�V�T,Ͱ�7	����'�\�2�����:5A��pfĉ>99��R�Q���~��p�������l��U5c��=�0��d������e�L �xc�e������C���ð��T�ݚ�Н�?V��j�c]���I���Z鎬�������(���kO��u�-%f_��m����ϏQ"j���b7�S
��n@V�� �9��1�Z���=���VvJ!�`�(i3�����!�`�(i3{k�h�+xއ5����-%f_��m����ϏQ"j���b7�S
��n@V�� �9��1�Z���=�-k�)$�>m�ڨ�hծ!�`�(i3�5ߧE4��!�`�(i3�5ߧE4��fĉ>99��A0ok�׹�����REJ���}�Z��/��;��|B>)p��I��Y�-?�?����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Â�	�ҔD����Me� 4�(�V��t�D%�}�+=&��:n��+G c��Fg�Y�:pR�'I4�u�������ea���Jm�W'�׏���15���{v���=RG�G� |n2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�Cn@_�b��Մ\�;+Ώ1;��5�}�]�����nv��~��i3�<iK�!�`�(i3��?��%��h�r�Bi�v�V���;AD�%�	-=N��ݚ�Н�Պq�Y�.��x���"x����O�r�1�B,X:!c*��!�`�(i3?!���l�~�y��(<�z4G-�vN��Dώ����ݚ�Н�Պq�Y�.��x���"x����O�r�1�B,X�굑��� q��j�J^2Y��kک����n|�p[Y���"�td���*:غ��4����ݚ�Н�Պq�Y�.��x���"x����O�g)�X��m����6 q��j�J^2Y��kک����n|�p[Y���"��/�`�����Y��ݚ�Н������L�	f퀔���἗jc��{��sۍ�s�*l�N*Cdr�3��15�\���'�s���C��E��R%E��g]ʧ�{I��	��JB�%OU�i�Ɩ��]�W\(���;AD�S�/xm����r�in��oK=��\I@�ZJM)����d�8��⺞=I߀%)���Y��fh����爮��J������L6�>P�2-i_m�;Y'�V!N�'�y�G