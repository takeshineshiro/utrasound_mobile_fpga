��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�����|"�L|�w.j��6��H4ي��2_)��:B!�b�ؐ:�{T�{df;���a,�|��4�Q��T�*0U1�1�:�Ω�����|"�L|�w.j��6��H4ٳ�k.w�.u���ŏ|{T%�at�3������ͧ� ?�ģ�ݶ�Us�JG�DGsc2�aB�>�;�C�l���o �����$[+r�bH7�D�C|N��^ �}w�*.��>��'��E����FDR��f��Us�'U�?K4��G%�L���om�Q*���T�K/ZT�@�t���@H���n�GE!���I0���������]]g�2�K���<�����*$��`�����$�^j��ʾ���g�����dK��m��sN7�H�t��%2�1����xZ��1d�n|s�)>��{����YF|q���#bdE7Hz�
g,UiB%C��g�� 6jy�u_`D�EcX1�ǝ�(�Z�6�hU�ڜ�����"`EQE�q��Ŭw:P� �����:uW��l�j#q���Bf�H>A��7`s� '�%�I��v$3Y��P4���d�*���%��38���E�!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�/�tw:g?�y��h�I����uk1i�f1?���b1�F��,��n�2��C�`Q�{���_��Bpш�#w��s8[Z�xZq��t�1�:�Ω�`<4}��o�r� ��J��ݪ���AOge���ئS��.V&��B֥+��@-�-'͏������y�g�M)ԉ���S��Lq�^]�+@���k��!�`�(i3��TG���PIÙ=�H�ܓ���A�.�hQ3'w�o�<m+r�X�<\�!�`�(i3��TG���PIÙ=�H�_�/��!�`�(i3!�`�(i3!�`�(i3!�`�(i3����Q���~������u�[��	��AɖD��L��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3@���-���x��Y� <~������'abW�5�}�]�������u��4];ˍH�7��_��T*�7⌹I�!�`�(i3!�`�(i3!�`�(i3!�`�(i3g�o�3���ء�Ch�1Ǥ �)�?�0��Y��W���ǣ©��!�`�(i3!�`�(i3!�`�(i3!�`�(i3c��|b�u:�]X��w�3Ɇ��C��ǟ�q
_0�>�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�q�����]��aT��0F��� }}�,���+�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i30d�N��H�ʤ�ܔn��aK7�������Ӧr�[�Z!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�aiM�`5�V��On�W�"�Ů7��B����;�K7���'n�^0o��~+�ݗ!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�S�'���� ����}`�/��+�!����/wފ����!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�|,��@��{��x����S����W�"�Ů7�6��,�;/�"���'n�^0o	uZ_�x��eX+��f�m�����;d� ���l��
$��3R�l��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�
ۼ����F#I�%�[<c�=, �	{��Y��
�iC!�`�(i3�����5	���]���>����C�Gظ0����!�`�(i3v�ј�"��Z鎬����F�71�B�������%�!�`�(i3c��Et��q���U�Ƣ�cP���:n##���Ψ�	�ǳ�6ϔO��)$�I��"�,�>E����-��%M�rs�i��s�٭���lC��U�T�\ ���A����_�Qf%u�!�`�(i3��(�
t��Y�{'%s�Ǹ2���;�¬pX��g��U-�eaԗ5��C��U��_D��.V&��B֥+��@-�-'͏���������6��w�>P�2-i_���F�� �yz��$6^�}� u��=��5W_�Q't�>K��cEp	���>P�2-i_��VzFI)�.�����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-����9���
�o�u�/(�,�A�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��n�g>!g��*��Q����aYM��_G2����4V�H�%�8I�_�ju:�]i�a�*��w+J����mw_�j��7޽.6}��bxUr�d�+�ĺ��Y �6Cγp
�얬Ϧ^c!�6c7/��.㟏��Z��/��T`��#�$ݵd;DuOw�!�}����g���ƒ���XpɽP��]�!��	Ǹ�y85��3}�@�7"j���b7|#9���\o�LCd��d5C[�[��蟔�,����}�쐑�8&���I|s�g*n{��7�4��~��~TX�'v�F��$ BŊ����c������ޏ����\�'C#/<���q���eacߦ/�;q
Db%#�'�{b�!�_b�ȅH*�#R�J�v��6�:�bt��l�+�7#��.`L+ކL�t��nЗ!v=iK%B�no��R]^�)��]'\gWg��	�Z�kfc��2���8���+�^n=\f�5>�|��ea��:�>�S��;�jmT�#bs��2[�a��o���zM#��m�!�`�(i3NL�Sfo�r��n�"��Wr���,(��9�e���}���|��p9�H�4BM�R'cf���}��Sa���D�#�e��*A&-�Ri9�O��F�I�؉P�=<�6>e��0�U+�qbp@�!�`�(i3fF�5.]����}Dq�f�����g�Z��3��a���!@�f")z.��W�����F�P�7��S����_�vL!�`�(i32�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pd����^���09���R��d`O��� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�ݚ�Н�:
��x�{�\��N�Ś�-����!�`�(i3B��C8�41����q+�=��Y�$����}Dq�f��V9_=(' ]���`,9�H�W�Ĕ���e4FgBĎ��Q?M8�f2!�`�(i3B��C8�4\��@�EB��C8�4�{D��ˬ�!�`�(i3�u��A�0���򴶽!HN��R��F F�E̠$f��_Ub��7��G_��$�)�vx|��ea���Ec��7�ꢤ�Og]���I���B��C8�4���2�cU�S}�3�U�.�g3Z�7�4��~��~TX���8I��2���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�+�DPy�#������Z�6�hU��/�����i�ڿ��5�Q��7h�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��6]@ÿ��$-:��!�`�(i3!�`�(i3;/�"���N�'�7)hCγp
��fH'��!�A���%��gx�n�޵$��æq��͵D�����R�p[Y���"�$L$E�͆����~�!U���4��)�Bi�v�V��2*Q=F��j#�{D�A�W+��W�� VU+I�A�+xĪ
*�)�v8W�����%kRq����!�`�(i3#B��F�!�`�(i3!�`�(i3�M>y
��;�?�կH�X:��+�S�9;/���!�`�(i3�E����F�׈PzO�e�n�^��$�)#��I��H��.��n��s����X=n/a�τ,�e>%�����!�Ȁ�k)H�=gq�!�`�(i3����u����\�vŜ�}Dq�f��am.�!�`�(i3!�`�(i3;/�"���G�Ա@\!�`�(i3�:5A��pj�.(Wx*!�`�(i3��gń�f !�`�(i3!�`�(i3��(�
t��Y�{'%s2�ew��5�%]���a(􆿳����^��3Lv	̅���8�u?��I!�`�(i3Y%T��BPe.��xu	�>��l%i�-��hy��jX�p!C+!�`�(i3�E����F��j��\w��0]��+�t2��ʄЀs�!�`�(i3"�,�>E���TD���rs�i�نW0��;�¬pX��g��U-�e�,���6+��V9_=('>3���T�!�`�(i3�����5	���]���c�A�L'�{&j����6��	�\�HP@�a!�`�(i3$r�t�}i	��D܂�Aeii�'��ƫ�G���@�|ųt�����n_�����S��ȍry��	.�n^y���\+��R�4.����P}ѪMjo�t ۦ� ~�p��ݚ�Н��L�K��%<7�`+Al��R��
�V_nu�$�F5k0B�#2\z���L�f�\c`���6	D�"�,�>E���	h��IB��`���oX:��+��b��v�#$�q�
k�E����F�׈PzO�e�n�^�(��.��dLG���6!�`�(i3����X=��}DD����}Dq�f�s���eZȗ�ET'z!�`�(i3;/�"���_�����ݚ�Н���*dy�ZB؋�Ly�H!�`�(i3�:ET֤vKN��B�)Y!�`�(i3%+bn/�{�.��8z�f������M>y
��;�?�կH��a�}�$Ϩ�;?���*/�|��E����F�׈PzO�e�n�^�
 ��4���>�*�!�`�(i3����X=��}DD���ݚ�Н��֠�������9���ݚ�Н�7�N�!�`�(i3!�`�(i3��|g�Y�'���Xw��}Dq�f�<9����!�`�(i3!�`�(i3v�ј�"��Z鎬����7.~t=� �^=^���3!�`�(i3!�`�(i3Yl���#�]�!��	Ǹ�y85�2�Ԡx��CyW�f�tR�wX��!�`�(i3~n���,a!�`�(i3!�`�(i3c��Et��q���U��ݚ�Н���퇇М1!�`�(i3!�`�(i3��|g�Y�'���Xwd�n]NْJם����"X��[�'i�!<�!�d�<HN��R��� VU+I�ԩ�V���5����`K����[���K�Ew*��XP��ȷgCu(o?CK������к��Y �6[\.�|���\_9ͫ��G//-���$��Xo�q	���߉�(���G
)w�<�_N�h(����.]̌[�$,��;�^P��:w'�>ſ��D�U�2Y�]�N��&�j��O" w��E����FZ鎬�������(���Jם����"X��[G�f�ȑe 4G�1����B�No\o�LCd腀J��R��e���b����+�J��Y�{'%s�Ǹ2���;�¬pX��g��U-�e6R��h�޳�������N�2߄�}�
�?�����湡N�Ւ>��4p��Q�
+\[$Q��
�̞��>���L��,0��Fb�E�[��Q[R�7}�
�?�⼲Y��pJ�V���Q]� _ό���.ӥ�n4s1�+��uK[F_Nr`e���7!ךv��� 펿��1��`�mp8V��0�$� ����9 ���Y �6���Eb�#i�@��՞�gx�n��\0��6W���k<��ЕS�#m,�?�d���&�������y�F_���ٱ'W�w��fD���ӽ~ZH���+���$ BŊ�J/u��xwm!z1��,��|g�S� ZH���+������wWi:rö1M(7������ȓM�Me��=4�pu��#O��+������.���!�`�H�� л��W�Ep�_���ޓ8���(�6k�4d��X��'"D���t�T��?E-h��$^(?��"��K�����+�^n=\f�5>����za���J�LQ��w�H����Qw�c4~Nr_�mS8<�n!�`�(i3�� л�4�>������9�@f���ʦ�/\<���tݻ�ݚ�Н���͝'�һ����e��0�U+�qbp@�!�`�(i3����g�Z��3��a���!@�f")z.��W��.�
9� ���(ٗ.;���JTv�䵪���l����� �'����u��r��!�`�(i3��o�	�=��Y�$����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t�Fr��jr��*�tzb*yX�ص}�	76�&�;��|B��vL�7&o���S}AǞkr��/� �~邔�f	�0�ߖ�P�T\hpo�h0�h�#"
s���
���b�Ի�!�`�(i3!�`�(i3!�`�(i3����"�	��J�6S�# [�T6��f�R��x����ycw��Έ��[i_1|`�L@�7�Д'��uW!�?�d���&�C#/<���qUI��������y1=����h�Y�X[�� �Ω��52+�F$0y�ׂ�G�3>q�OG����SM0.�,��ʇf�c|���p���rJ4{Yp o��`��:*������ɢX��4tΘ���=+XRw�a��$?�C#/<���q�`Ҧ�׶�>��Z?2G�j�W�������o�u�/"<)�]mY>��XS�2p�$�����KCgB0�/B�xiI9�o�?�d���&�3���L=l���ӽ~ZH���+��M+���C��v{��lw	�m��^�����,�ǰ ����U��X�l"��h"�+�r���)`s﫱Och�����ƛ�������l�`!�`�(i3!�`�(i3!�`�(i31M<���8�W�"�Ů7��B������z>9�R��d���!iO.C�+��uK[F���Aw9����Och�����ƛ���Id�U�mu��0\� ��+2a�u�=�d�tar+J�Y.i�t�cx����y�mZH֫&�9|�CL�qߦz#�� ���HoF�g���A��̙(^���/�RvE�3HN��R��?�d���&��n5����=�r���Q�H����S
��>ߓ�~��O�1�l��g@bong��*!�`�(i3!�`�(i3!�`�(i3Y%T��BP��Vl�8b�m�N^����d���!iO.C�+��uK[F���Aw9����Och�����ƛ���Id�U�mu��0\� ��+2a�u�=�d�tar+J���C��bU�T�4��uZ(��4�WT�e!���1�~w���?���#�"��\�fh������bB�o?\�z?Xk�V��	��yAsr�7���X�u��ȋ�=�^�Ne�M� N&$Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �k�����f��v�����;g�"���	�VH�/7�4P)Ɠ[v�Bx!B.��(lD�������<�d�:O���@B�d�G��ݫ������Z��r%Ʀp����y1=��_U0�H�/7�4P)&.�P4XEh1�MY���%��u��p��ν(C�X��4tΘ1�E�Ou��"�*���h]�ǚу��+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}ژ�O�q�:��&�̎!7����[�2�G�<K���Z��C>��Ӛ|s�g*n{��j5�{��j��(u��F{/���s2F\�M�jL��Tt���a lϗ¾IŌLNk�#������%kR��������֢&@��&X:��+�<6��$)K�X;p`�#B��F�f�?ǉ�=(��.��dLG���6rQ�4��+�I�P�,���-�X�fw!�`�(i3*�n�6��.7x4�"����5�q	�!�`�(i3D��)�a\_�@ ��G
�/{��(Hg�"�I��6��w��'�k�f-���
�I�>y�ݚ�Н�������s�e����kn4@Q�/�!�`�(i3\!{<�NM|!�`�(i3�Fv,"�_O�[��?���hy��jX�p!C+�X;p`�(����鹁+�t2�,E)�ک�-��f6ȫ�-��ݚ�Н�k�k�c7!�`�(i3��{��W�mOeTky�!�`�(i3"���
w�&8�,��#0_K�>!�`�(i3�֠��������,�ǰ'�J:��XD�v*G��tt�td���5�p���C�S�&�̎!7����[��t
����Z��C>��Ӛ|s�g*n{�B�ek�5W&����]�¿��L�j�=D��W�/�#+*f��s�vV�!�`�(i3���^���M�_"�]*Ò��u� ����,�ǰTm�v��G��G-"ұ��5݈��]Ճ�������_��Tq�'?_:[v� 5 x����ycw��Έ�͌��t�h��W+��W�{y����M�V<�'���v��|�>�B���m<�6�Q=Pip<ɯ�n�^�,l.8��J��G��#&�Y<�6�Q=����ըi��D�].2���g�ecVu�RV��,����>�v�䩲$��߭�?8�)(����<m9�����5��4�Wq�2�QR�e��zԶf~���\����6�o8:4�I���c�90�Ǘa��x[�����:Fa�7����os�鮊�� ��9ڞ
i�c�r�xjzӝ���I(͂�'�ɳ��!�`�(i3��4h�=Iz~r��V�n��dK�����fF0��!�`�(i3@ E����/ ���we��0�U+�qbp@�!�`�(i3����g�Z��3��a���!@�f")z.��W��.�
9� ���(ٗ.;���JTv�䵪���l����� �'����u��r��!�`�(i3L�,k�6�"%�iq���l[�Ƶ�1tSjv�!�`�(i3{k�h�+!���?t��my$�N��o�/���;!�`�(i3��w�w:�!�`�(i3�2��}��e�g��)$�j�=D�Ȝ�}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ�U`������kLZ�.�g3Zdj�t����Қ�"<T���Y�b��K��*� n2ϒ��xi��?P�dݯ����o=�Ϧ^c!�6#!��׏��Z��C>��Ӛ|s�g*n{�Cy;"-�>�@��<g$
�1d�9���c�}�p�n��W�/�#+*f�P~I��ñ⼲Y��pJ�V�F!��D�����k$ !�`�(i3k��_� ��(ӈ���m�r����w�R���yǿ)~L��"*N*�i>_��Tq�'?�Y^y�*ܦ�s�m�d�tAgo�\�<
|T�!�`�(i3!�`�(i3!�`�(i3Y%T��BP� ����9 �K��2WI��z>9�R��d���!iO.C�+��uK[F���Aw9����Och�����ƛ���פ]�|N�C�7�/�)hΜԹ�f퀔����:��4�_�2*Q=F���q/���<�9|�CL�qߦz#�� ���HoF�g���A��̙(^���/�RvE�3HN��R��?�d���&��n5����=�r��"�U���50��L�r:Pip<ɯ�n�j(�X-��+��5K�����s�#��OƜ'�D�m@/�%�\��l�]�12Y�H���3���O�Cԕ�)>g�k�4.��>���c���v~��6
�@{>���q��M�$�F5�YY�ʙ��9��ݔ\�Ϊ��:�B*�2���h�8l���>&� �V$Y�4Eb���I!����)��Uza?�?#�*�bP=4�pu��#O��+����UD�5���c^���H�k;��7O�Z#br�:l[[Oթ�߁��8�E�"0f���U!#����"?��A$�P������5d�`UNP�{y����i�q,?5q��/�TPe�[Oթ�߁��|#HK��A(�c���_G��Hb�8�u?��I!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"�4���i&X��7��C�lԇ�-{ÎD9��ɰ���|e"/w1z��ӊ#���ꪆ��Lt�2�tE�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�7<(�lb��� л��E�BS�+��U�,�P!6���r�����$XR�QܛOcOZail������&G!�`�(i3�LĻ�ڱ�Zo��?�{g����L��,0�tH���b!�`�(i3/w1z��ӊ#���ꪆ�'�������xSC��k���4�b��~$�!�`�(i3@�=�{��5%�iq����/���bx���NM���
�:qEp'{w#/ B!�`�(i3&�H
�D�h�����0��$�\%e��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��/�TPe����z���;_��8W�w��fDy+�gr��w�1N�&�_2��VU(��z�j�Aa�R�