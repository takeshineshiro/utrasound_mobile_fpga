��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR���b�z�>}��������M7\F���r����&$9g8�M>PFWD#�z":���ӳ��_}��0w�\��8׋�������N���?��m��+�ڔ�wV���C�Sy6ג��̹��/R$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us��n��/�FI���O8�yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��7��ri�Z�#ʹb�r�	j���@N1�w�0XL���t�ے����o��f?��n;�|-���g]�܁��U?���S����]�jz�Cb��X?B�/�a�{���r�hr�W�M:]�Idr����&UVa�(��z�j�T�٥��Tּ���)���C�\�T���WӕC��D��)0����,��.tK�z':�
續:�5��f�
!|w�̺f|��/���P�΃��V�/��=c���X��d��9��G����a�����(�I�?g�f��m���b�� \
��툑E�TJ	V�+�N<��;���u��w)�S �J���vy��e��m*q;�K?���p��O��Of�+���jv���z-&)�SD�:�Ä�����N�v����
��e��o����1�����(��^	�܍�1s��i.o�*nŐ�u�l��êME���W͉A�?����i��vp�$_<n�ȳ؜k`��Z��L�R�.�$m>�-�_]�og�]�n������fxQ��)��\�4�s�gD�bOq������ǃ�8ƶf�,w9������ֹY���8C�j:`d!��tW��] ��[+�c�5���AQ� ��_�^�r]��K�X��K�zb$z{
� �AH��T���x�3�Z�<uo��0]��;�*tD�>;�L����� ���>	I�멲ٰ�Ř�h^������*����	~+�<���p2��O�_Kc�[_H|�eĕo��tW��] ����&�[>�y��W�y��MqZb�L� �k�#�l�w|ü��}T��X����::R�nҎ� ��k��_֦�j0V5����
� �AH�h	_�fx���Z�<uoz�!Կn��i}3�L����¸
uy�BU��f%%eo���sp%S�y,Y/�7{'3'�`�m�!=�y����h�}K?c�*�S�\�l#�+ohCoǬ��oB;sѱE�?�m��l�j���N�=�����q*\�9X�����XQDi����N�v��<���P���d1���P��)2R��DU�AP�nJ���_U�t:�W�g����J%�hu}�fO`�|�2z�R��톋%$ n��c_�Jh�5L��p
� �AH�+�6�O�_M��RwM�麶V$�(k��n�L�����r���(�����5ʦ�&�d�I�_ K.u0�p���?�o�3�P2G�e��-�u��w)�SU��T�d�I�� ���I�"{��&U6g���Kf�+����Z��r��p��>����}�F��qt4$p�)�����W{��!�*��x�6p.��k�8���҆�|n��tCP��뚽���I;������4I�0��U�)�(27�׳������<�6�+r
�M95��v�7����}ʬd�ŷ|�v������s��"q�Aj��6�T-t���S�X��Z�Ʒa�o�u�/�|?F���DB�T���xĄ}R���~�$�Z��ДJ��_��"SӠ�|&�:h��_���&Y��V�F��2��+��T����5yi���FnBƕH�N�4�TLAZ�Mg(�}���Gj0�0�G��O�2ҙ(�r�O��C��0��/Ί�lz�NC�5�+D�)4Z�|p������]��b�4V�U��}VsTq>9+�d����k*�Q����uc���&������D��������K����J��\�4�s�l,�(~�Z�o/5�i!����� -hp�74<ֹY���8���+��"B�A��dR��Wk$��X�~�b]R�U�W�M��m�!=�y����h�}�k�{w~2��Z)H+�`�Z����oB;sѱE�DK�\�h����BPMF�I0(g>�90W2f��j�]�}��:�����,�A-���:=��|��۱��@5Y@�,���������\�4�s+£>�,cMZ�o/5���#h�o�jR}_�ֹY���8�B�(�}턋���\��>��+�q�������c� S,?[
� �AH���ಆq��M��RwM��P�	�����~&[#a�i�L�����\n����r?��,��T�X�P@$ �l�q��M��ew2�\�����	x]�Ħ1��&�8���X4�c���*����|my9�S�O1���_U�C�s� �[�|%�-���:=��h�7��sB�|7`��w��RL�a)H��dd�@=�~篟|�CY�y��`2�-9�$9����E�9����\`􊩦R�L�1���Ajn����p��8�hHh�<LXn�r�O��C��0��qY$�!�",nDi��
�V�Z,��G"�C�"���<<���E�qt4$p���tZSA`m�!=�y����h�}cg�I��O5|�iiG�&�/�b�x��oB;sѱEϼ����=�>c,�©(��g��b��S�aa��2��9�;P�@�S�c�@�m
� �AH���2\�����(�Y���mT����ʋ8���r	�w�L�����8���п�ߜ�I�	U�m�!=�y����h�}�
"�k�'ވ��#:J����)�:�-oB;sѱE�v������I"� �����\~K�f�h�9LC=���\�c[b���M�X����>5����A=/m���9H�Z�ǵU�{�u��w)�S��X3��¯(^k{3��R�!�"s� ���z�?f�+���zI\S7�8���
9��HB8�	S4�"-huڦ�W�PEQQ��ƴ���(��}���W��n���3�=ذ{	���7ߩ�k�,��bҢz�n�j{	�	m�!=�y����h�}`29�$zFq�Be�y�P�;c�95oB;sѱE�'�?��M��N���p�U7�"%��-=���"�9 \�/�!���k�8���҆�|n������A�"�K��l�@�'"ǿ�:�����NS�O1��Dtr�$�{���R�������	x]��>��M�}K��l��A���P"�a��R�S�O1��{OE�c´M����R��_��4zV�Ė����D�P��w��R�k�8���҆�|n��Ϣ
[FH��%�KS���$�Q������U�)�>(��m���z�#˭䱾n}?C+�׆��T�uXSr���K�d�eM�bm���� O������C�(#����{�;¬>P�2-i_)[���G�N�Er��oIIB���?��6�
��G�܌Y<����O�?�1ag��vu��w)�S��X3�����@��."�1���o=a��O�f�+��������l�����~�W� ���>w���M���o�G�m�?�蜤ޝء�=t���\���*����U��+�Xa�H(�˕��as^+�t�k�8���҆�|n����:Vx�p*��&�BSz�q��f�+���X�LGA���oS����Bu�����	���C,�o+P���f��y:��c��.W9�5��H����-QpK2'ōeʣ͜�������t�rK�gRL���7T�y3�Ɔ ����uvo�N�Y��Xo���1B�:ͫ� yԶo���\�4�sƐ�hd	���(�Y���m��V��J���	�E���L���� �G9�lF$����ٗ���吓z�>��lǐp�~ZQ_%8$�0/�� m�!=�y����h�}��b�Z�ԃ7��L�(��$�'z���U�)���IU��_U �mɗg�T�~,v�H�UJ�r�O��C��0���۞�^�(<ڨz���wÒF�oB;sѱEώI�ݝ�~N�o�L�����RL�a)�ƞ��U<�K+8�M�����T�%��Na�ֹY���8'U��&�f.����S����?�~����\�4�s���rH
>�(�Y���m�** ,�O&��3���L�������"������l&�ǿ������F�k�8���҆�|n����e��m*�R���O��kή�f�+���`��Vԯ?� .���9��3��F#w���9��d$Ǵ���G�����m��d�7��v�5ܗu��f��̽?�4�ʗ��Z#�!,J�l�/a;����XVx)ۭ���,��m�Qp��)��	��a�u�$f����D���i����	x]̍��;���9�n��j�ih�3�T87s�!��O�e�'}�����Z�4]u�t:�E����jp���\�4�s��{��]Q�X �9W$%��y*�vc+�^\L����� ���z˞w$����/y!Z�5����5�"�IN�RV��'�͉�VZ�����XO8��/�:Y� Y�@����L���W y�!OP�n'm�2e�+>԰�A^T�?qI���"����Wv�A��xİ k�����
r$k��{0��d#h���o4�e^�G��J[�f0� ��[	�V���������7�:_���.��51��SK���B��翑��HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A����2�P`��������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc$��+�{c"G�ۄ��O���azhݪm����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s��e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3����M�	g�y�+��T��C�NJ���1�:�Ω�A��>s>;����Ms�JFAa��Bzb;ym��+r��JʅY�y��
r�(����5�����x%~Y�1�:�Ω��
�/�rD���J7"���`���lY�y��
r�(����5�����x%~Y�1�:�Ω�S�T�;Ϗk[�^��_E$ô&y�#�̔"v�lf)@̲#;���(�s�-���f�i\􁗊�n��\v;V[���b�/ri�y�!�3]o��in�m��+�ڔ�wV���C�Sy6ג��̹��/R����h��,��B	�^�e��I�	5��2�$���w'gx�r�ľ�q�ܺv7M?\���#�^!��z��TJ�q��r�[H�l׬o-ӕ��J�U�} {�m�����`0r)&�1c.�Mn�4ҹXH�A( ����_ֲ��mŹ�ΕA��l�='��:sF��Thw���иܖ��i (LW4�'n�^0o��g_'+���ԏ�4��I7��-5��;ε��IÙ=�H<z,Ҽ&�כ��p�k�c��`��'n�^0op40�zɈ���y�,@���k��JHn��z�:3�>�<5��Q�[TّD ����R�^Ƒ���b9����4�6�t��e�I���&���5@���Ml���Q**�7`����M�Z���	�b9����t�V�h� ��S�����B7�B����{�����N����e!M^С$��JHn��z�Sp�}�f܀�(nԐJ*�Rs�08�b(���b9����pP�o��a��cn��;���N�H}ة2�IÙ=�H�M�U�h�5,Wlr�r%)cA��u*K6HT�����N��2�F�P��U��+�Xa�H(�˕��u*K6HT�����N.��TQ:-�"E&��� �
�V[�}rYs�7��M���HaU$kX��� nU�IÙ=�HF���m¡A�h��+Fen����9��#�B�sYC��\�v��_�R�G�$����{v��G�K$xE�p4rqG7��u*K6H �i7�sp>��%��H��5[�����q�_�N�6�Ặ��Ϊ�Q� ~�����(��q�
�Bk�i�E?�xu����ma��u��ۯi\�q���Ì �&�k��>���c��d�|ݔ�3�5�}�]���x�]�V�����Ү��`�+S�p��ͷQ�X�����d�� ӫ/��m�A0`��A��L�>�c'�'n�^0oa�䪱R�JI��_��3�.���˴w�T:~�b9����4�6�t�P�(��܃�mD�o���B)|D��P�Sb�^{?	�c;5�}�]���x�]�V��7��_��T*�7⌹I�Bg&��C��5�}�]���x�]�V��7��_��T*�7⌹I�a�ɼ�Ǟ�7�/�B*�7�ܥ��2�)gvF伉� ɧ)�2�X�S[BYI�kU��94˯e�B������.�)�p�gR� �ұ7�ܥ��2�j*؂�5�����\���a
��|���\G�Y����-�,��Lt�2�tN�By3��<�]�!����M[��Ǣk/�z�xEQ�����5	���]���>����C���"����Y%T��BPe.��xu	�>��l%i�-\1��pz��S⏸[��c��Et�Y�{'%s�h�v���5���T�`�|��K�z�L;Л��Z�n��[��{_8�Y��=�}�Vݨ��������P���Qi�]2�y�Z鎬�����,�q�����CsYl���#�]�!����M[��Ǣr�x�e�X�����5	���]���c�A�L'��!�a��5�%]���a(􆿳����^��~�ӵ(r7H/t��)��-��%M�:2QYeƈ����OǍ�3�f�P�o��h�Xޓ$���]׽������E��@IE�U����S8����;(���5�%]���a(􆿳����^���#}�{�,�k,^+a�@IE�U����S8��$FW �9�װ?�p���5�%]���a(􆿳�ؖ��d�I�� �:&��I�?g�f��m���b�� \
��툑E�TJ	V�+�������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��q�©��7��#!l'����z��d��o�vC��9���$1mT���u�I�	nrB��ZaԘ�������յ�}$|~ïSup�xg쬉� }���n4s1��7�癆cg�!������:"�9ʮU:���s:��t�5i^��EQ73)yn�w�x'���Ě���aT��3G��?�#M'���"��y��6��S3�ߟ{����c�,�V(��_�8)$���}6<6zY~G��A( ����_ $}��}5Xx�	�+�&I(&�L�ӵ��)���>�ѻ�5����g����ĳ��2S����"ܲ�����^Lma��C�<�Sm��q��Gh�3�!1�F$f��_Ub���uQL+����6��S3�ߟ{����h~E��+m���L����Ҙ$7o4 l�5Y�0`�WC����B{�LϬM��+��!WS���
9Wp��� gؓ��')-W`������a�"�fE~�cb�i0[����8|��`��W�U	EX͇�jO���a��Ó=�vzFg>"�vA��K1P��)�b���g��� ��"�~�>����;�P�t�5qM�4��o�Lѯ����Qٯ�b���L����Ҙ$7U2�h=c�ugÕ�KF:����Į��KH ����p4c�.�U	aw����Ѹ��ln�~8!��vp�o�6��aH7luP7���8-|�DF
�j��6������1�R+-h]�0�tW	�pg^��Pv�
�\� �jO���a��E�' �!��"� +}Z�"��%o�&��cay�[}�	76�&�� Ӗ�t�t��"^��#��Q���@��q�r����開s��m�z����9C��,ў1�ˏ�~ǹ�z��hbvk~�#x���EE��n��V����#���F�O��$�}$|~�﫞��fS�Q�S�T�=k�Rm��̍$�D�u&g()��ikp���H����-��԰�3�#���F<�X��j������&<v�}����1`�O�t_)x�?{��J�SqVEG��5���-�;���N��}�!`�������a�"�2�ʏ�"�<��E��b���a.Y�wg������F��O�z��K	pgu�5T��$ VRMR��,�*�K0Wi�l�U����;�� ��-�3��&Oa9Y֪{���ɖ?��_T���a�aq��ڷF����/woP}[�.ᬵy��5_
� �����3���ne
���HK�0,���U<� N��r*�jB�B[�)x�?{��J�SqVE
7�Ԗ�E�.ᬵy��5�H����;���<@�� Suiӑ�xGe�;���N��}�!`�������a�"�2�ʏ�"�<��E��b���a.Y�wg������F��O�z��K	p����)Pg�ŉ�u��M�B��{���"���@
H$��j�>���?���B��Ul�~ǹ�z��hbvk~�#x���EE��n��V����#���F�O��$�}$|~ïSup�xg쬉� }�=k�Rm���ӑ�xGe�;���N��}�!`���Nj�a=�t[a_�?��J*�Rs�0c�툼��#���F��3�k�n�V*ڎ�0���J�և3
�v�v-}�	mp=b�ɝ:�3GV���J�1���-�".Q����>���?���B��Ul9��f;���"��y2�LpOJEl��Q�P�]zm?9ۄ��d1$�Q�<om���b9���M��A���va�{����U ��z�!e���im�th�U�CLB�D5�O�X��WG ���y�9�3��4��A�(bGuj}��8�,ԱvD3n�x(�i��/Rz��K	p��ay�Ȇ^���x�k]m���C�MV���%��b����3X����a�x��M�ݭ�~r}*И��&�������Ŏ{�"��}�偢��%�<ͯ�G��R'),��`�@ux�[����3���ne66�v��G���V>�R< N��r*��حFہ֥��ع��8�b�R$�Տ���i���a<�*^e��J�v�t��Ʊ�_�eD�I��3��oE���$�8@�ɮ��U���#Â��&?��Nj�a=�x^1⩠�^!�<8qx(�i��/Rj���;��D3X����a�x��M�ݭ�~r}�֫��XA��Gm�o�j��`KL[�{W�g���F�i;�:U�v�3b��{"���,���"��y�xI�2^)b��@ŋ��5k.'C���Y�V������p�0ty�P���Պ�`^��3�J��\�v�w�?�b�>޼�\�vř9���=��\���.@A�-�]s�(_�<�� ��b�FP&����҅JHn��z���������x�&�F�]:��='����R��e%�2�ͼ���y�]�F�D�+�:�G�9�E᭗��_��&Yd&�j}!��n�͑��LK.I�:���3k��g1�e%�2����莇����_����~���i�x˗9��6�8�d^�ϓ��ͬz�Ť��xI�2^)b��@ŋ��5_@&:������;�R�I͗� �-�`)��\^�#�f�R�I0���ԏc�r�(���JHn��z��|/��N��hk��Y��A�m�(�b9�����閝eu�m&� JHn��z�w�<¯�����v�8:®xԜ��H1Y�ΊS&h�5,Wl�/�O'�=�ƣD��8!��vp�P}��O��^��mi9Ů���z�jaV�,�&{�zYa䃾���Kl0��F��j!-`���w�|ò���
��_��������[a�[�J���6�@3uå��:(�
�*S�#���F)�S������4���XP��ȭb��v݋N������5R܅dJ�A���ۖT��Go1z�Ů���z������e���ݟ���O�͛PA,qLn��S�W�
����uK�r�&U������G|M��M�~}�]�+U�HJ�h<��}@�ͫ���r�3�����!%Ah�%4
>�(_�<�� ��b�FP&��獶���_�(�X�)�v�V�.��b9���.M�"��Ӗ��s��2b���!h�b�TG|�w57�S��pN��B�)Y�+U�HJ�hn�./�������|I1=��%Ah�%4
>�(_�<�� ��b�FP&F�W�1'����
3��FZ�ޑǇ_���˱���v�0���f70���!�`�(i3�����5	��M�-��#�g#���I}��NV�MO���9�<�!8	�I]��� N��r*�$��ûX��kRCլ�����`��&f��w�'�?t�kJ �&{�zYa���<��ɢ�U8��ّ�k���H��@!�#-�[ҭ�g���y��b��v݋N��������c��>z�Vg.N�������6���|��"5�o٥۪	�}a�iQ��ׇJ�	�LÆ��/�i�����܍w�S}9g	���W���b���p��=�^���3
�v�v-}�	mp�����2x�N?Dd�-$#�0$�.�-v�Μ(4���Yk˃Tc�δ�0���'?Rg�\�G���nQ�rV���1���X��WG ��D����jF��b�(� �	T�����3
�v�v-}�	mp�cA�N�Y�74��LM�(�� 	l��lBýO����ezꥦ��r���:�����C��괽���5%�"|R��9%2�8���x�Y�1G�Sזi�)x�?{����ҳ�ET��o*|�[3�^�P�qjhbvk~�#xe�����t���3��Μ(4��fU��S��ɻ�7��M����v�l5��� rư1�l�_�4��׏�����M\]YD�^�O�<om��Ts��E=�!�Wƞ$�FA��mӡ���<K�yw���-�3
�v�v-}�	mp�^5��$�9_��i�D�,����3�<�:@�@��\l�垹Y8��#�8���w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�w��AW�Z�y��l�Ow0H��G��9%2�8�Κ���@>��nQ�rV�����J [ܰ1��?�shbvk~�#x=�;����b��v݋N�������0'n�ڹ� ��yo�}�Y�PX�)��s����A���cZx�.��8wCc ,P��#��\��v�8:��MWU�?
�5ߧE4����{�A��3D�� <(rK�� ����ޙ���9%2�8�μq�T�<������t����==�x�Y�����5O�r�����Tb΃l�����}0x�PI��e��&�'��;���N��6H*��l�A���ۖ!���6�,N|��|(F9%2�8�Α��H����ָ������%N�ݚ������	5sJ�J�	�LÆ��W��C�܍w�S}&��|�7���Ɵ$v}�S滑���f�� ����p��}��aq���g0����Xjۙ�)��s���#Â��&?���J��6>�2�q�]��x`��:�x(�i��/R1`�O�t_)x�?{��J�SqVE�e�H:�I0���ԏ����[���Bf��0���f������C;�,]�eT�n
V~$�H�*x����=��:�H�*x��1d�ެپP۪	�}a�l0� �A(�i�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��n
V~$�Y���� ��@s'R�r���t;\`�r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�ܿE�qqRmF܂d�ۤ�m�>!��bT�$&�fe�X����)ͶG�q�5�
p��r%̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-���Y���� ��@s'R�r���t;\`�r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�ܿE�qqRmF܂d�ۤ�m�>!�����4c��X����)ͶG�q�5�=��ﯭk̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-���Y���� ��@s'R��E=���r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^��o�������|I~�I����uY�0��f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#L�tD:��@F�W�1'����
3��~�/:���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��'#���n�{�X����)ͶG�q�5�	`�/��í��H��@!�#-�[ҭ�nɦ4��De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�O�β\�{!ˎ]":V���"^Be��Dc]�`6X��3
�v�v-}�	mpҭ���^���b��v݋N��������;B�鉞(Q��;��b�=��?njS��}�vo;��|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*��'�/7Ii�^�Ax񣘂D-\`��EW+GE�Kf
�f�3
�v�v-}�	mp˜�ķ_�L�b��v݋N�����6�pnWwщ�(Q��;��b�=�`��N�G�g�r �����=}'t<��ġ��,.R��д=|��(Q��;��b�=���N��/*�A���ۖ�ꉴ�dyi#nĖ�*i�^�Ax񣘂D-\`�����SVc�Kf
�f�3
�v�v-}�	mp˜�ķ_�L�b��v݋N�����6�pnWwщ�(Q��;��b�=�
22x`8y8�g�r �����=}'t<��ġ��,.R��д=|��(Q��;��b�=澖f���e��A���ۖC=4�a,�n
V~$�Y���� ��@s'R�r���t;\`B�R���>_���!&�+��h�G6SX��Xjۙ�)��s���'��m�xl��(Q��;��b�=�ύ<Z=�	��U=��G>EK�� ��Ut�\��Y���� ��@s'R�t��&� ��"L?���J4[���w�����1��r�.Gb�TG|�w�q-2�;�"�2�q�]��7�H5�RF܂d�ۤ�|��F��ڊͣ�:Y��Y�^�f�s�tG�ه� �4�<��U=��G>EK�� ��Ut�\��D$��:��
3�t%9��&����1�%d6c�d	�Ȟ���p�o�QM�W?#<b��>
rw�&�z<aSm�6��`4�04�jfh�x#�L_����	�r��9��o���>6�P��%,��7n������A�9�-���Y�f,�s��Zrt�\0�{�q֣���óM�˄NKYi����L;ø\����?v���=!ߎ�΂l��=5;�D|�[�R�n��V���|ò���
��_�����,fF�7�1Y�ΊS&���0i���7����NT�<�*�!g()��ikp���H����b9���ʵ\���Ex�y�Zgl�[��j/Ҥd�X�VM�����a�"�'n�^0o.�ؙ�b�Ӧ��9���I5�4`UV#-�[ҭ���~����'n�^0o��N:�@?u�hk��Y��A�m�(xE8�ELE��&ċ�;���.{2Y��{�3�P���ġ��,�Q7I�2)��\�v�#�1�N�_�n�To�[��8-��-�3
�v�v-}�	mp��T�����,�v����f������C;��S���'n�^0o4��t-s�e�J�Pn\�H�4I�B�������y�r��VYW\�o���*ٝ�/�K^b�;��	+����4���XP���3Zk�E��% ��q ���h�c�M���v�8:mvvb��_�.ᬵy���=t/��g#������a2����b�������<X�l0��F��j�?��;
V�;���EWrN|��|(F9%2�8�������JHn��z��o�RO�v0I��'��_�(�X�w���vc�f70���JHn��z�9�Wz��
)x�?{����ҳ�ET��o*|�[3�^�P�qjhbvk~�#xe�����t���3��Μ(4��fU��S��ɻ�7��M����v�l5��� rư1o8�<����;���EWr��$�J݃����t����FZ�ޑǇ_����'W�=�-��/�D�ؒ��"��KH����t��(�z�=�j��\�v�Џ�I��$��cn��>��u��j�E��*�j�H��b�(� xܟ�,3JWA�%��fOX�����̏we ��g������%ng ���3�ҺIÙ=�HM�f�<�O���L��^�
h�tG�b��v݋N��������2����hk��Y��A�m�(�{`x��%5[��	=g()��ikp���H����zY�l��R�}vJ^��l�|- ��b�FP&�q���3B��*w�o9@g^�J<�b9���.M�"��ӖEKM�yW�T�s Wd2U����v�
����4��(_�<�� ��b�FP&f�%A�)!�`�(i3!�`�(i3�b9���.M�"��Ӗ����������
�x�w�������������� �1x�itLd�r:ha3B��*w�C&�5,���a	!33֬�lPCrM�Zc��~�/:��ǆQV���Ҥ�������|I�W����x�A/�n6�r\�H��/Sg4�y�)@��]��0�ȍ�x�>c�K����&&\�0���eYk�	�yOx(�i��/R�Ȟ3I	��.ᬵy��H *4�ڮ���Bư��9%2�8���x�Y�+���]���J*�Rs�0u����x/��'�ĮpYÕLM�(�� 	l��lB���U%�p�zꥦ���i͑��Ԣ���C��괽���5��g����;���N��-Lk���ޟy�K����t����==�x�Yu�~����J*�Rs�0u����x/�'��ޙ4!ֱk���p�˳c��sCF��[ S��x�%�/�d�"�hm�^�6/
��VLM�ǩ��8���׷y�S}m� 2�k#ʘ4��\��sپ#�J��v�8:I�}-��^R��	�ݑg()��ikp���H���ʤ4���aHUv�׿e\V��/��x�%�B���vs.�^�6/
ڌ����S�|���#q��iQ��ׇJ�	�LÆ��/�i�����܍w�S}���d����_�(�X�<�q��Dp��3
�v�v-}�	mphpL��m�d������g()��ikp���H����-��԰�3�I))����A�m�(ą���P4�=KmS��3D�� <(rK�� ���$!��8f�� ��}���x�A���ۖ��P4�{!� ��3�F��Zr�Z��T۳�͕��w0H��G��9%2�8��!����&@��(+���<om��k%-uב8)x�?{��偗#���\ԍE��C��>CR`�y1��r�.Gb�TG|�wA�2)q��FA��mӡ���<K�I3����b���z�òr0y4{�H�a�\�#���Fq������n
V~$�H�*x����=��:nQ�rV�)�YBa�g()��ikp���H���x��3�Y�^��q,u;�B�R���>_�qЕak֕��A�\>W�/Z�������u�`��3+��f������C;k�k�)%|�	�Ȟ�����hLKWX��WG ���
�����w��r|��߇(���л���.Ȃb�����V�I�e!��nH�W���:0>��� Q��!$�2�q�]��wc�}�![B�R���>_�?Iߕ��1ҙt&H����y�]x(�i��/Rh�x#�L_�h�:��p�3
�v�v-}�	mpҭ���^���b��v݋N�����6�pnWw���z3�:��c��%2���ʏ!�܍w�S}&��|�7���Ɵ$v}ֱl�40ߏ3��#Y�r/��5Տ4�04�jfN��������KG�5�zU��آ99BI|�6|����J%�hu��y�c�i������b?�*����f�����"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�t�%�(^?�f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#�P9(�bC�3
�v�v-}�	mpҭ���^���b��v݋N��������;B����z3�:��c��%2���ʏ!&f��w�'Xv��@�E��`;�nQ�ǅ�a�
ȍ�F�]	
~ao.\C�k����|�i�^�Ax�6�װ���='Ӏ�d&��(Q��;��b�=�OcDb==�7��%��Gy�ˆn����N��+�?ݨ���#2y�Z���7�A�6x��iY�g��ѵ�"xC��-�T(u	M^)FU9����g,Z�fg�4���R��T��̪mMUt��!b�4=y�(ͻ� ���7���ìL��-)6�oȔ�T�͒�H��@!�#-�[ҭ��:�*�3������w2}�<��bd?�&���u�~A4z��4^i�u�J*�Rs�0�|�:���@�����\�H��/Sg� c�Z�q��uY�0��f������C;�,]�eT٠�Y�����|O�\�+�q�� 6x�@�޵B�
�#�g�r ������w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x������|O�\�+�q�� 6x�@TW1R�X�L�tD:��@|��������2���t�I�� "\�H��/Sghg�R~G�����A��%,��7n��̥��}20����9��F܂d�ۤ�����ms3M��o(ͻ� ���7���ì\��2l����Q�=ؗ���`;�nQ��A@��sZ��o���*ٝ�/�K^b�;��	+�/��~�;1֬�lPCrM�Zc��ʪ<4 �"j|�S�
���N�@E�V)�jP|B�1��6�G۽^�w�򪥃�n�{��l[hbvk~�#xM+)�C%�&|���BY��l��=5;�B�8��\]s������&{�zYa�k�f}�Ɔ������g����;���NC")t[p��]s������&{�zYa�f���%��)x�?{��
0#`�1��n
V~$|��������2���t9�'��_�K�z��d>Q���G&o6��~��<o��!h�b�TG|�w�q-2�;�"�2�q�]�>��O˻����|I�w�63xHl��7=�[G��"xC��-�T(u	M^��|A�IU���b���"~6���aq���7��Y^&��fx'v�ao.\C�k�4yn����q���3B��*w�������(�Ae�̃B���K�<om���м�1#���q���3B��*w� eY�NA�J*�Rs�0$�9͹)��X��WG ������*��P3�lWD�q�5�=ڭ��"xC��-�T(u	M^ �(팵���$�J݃����t����
0�@lJ*�Rs�0K=X���d��h�e��SV�Cagi�"��(Q��;��b�=�U3{����B|�S�
���N�@E�V)�jP|B�1	S�%̌��n|�
H&b_�n�To�[��g���a��>�8-�ށ���
3�E�ʫj�>��O˻����|I����ZqM����
��\�H��/Sg�zH^x���r���3墚�w�ǻ��v�8:1~��vA�~�㕜��z ӫ/��m�tU0�x�^܊@3+'�tL�a.l�n�)^��o�������|Iܲ��9m����͵De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�X������<�N�����K����������\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���Г�D�i�^�Ax�`Vk���|�zYק�̒�H��@!�#-�[ҭ��F6q,/̛uBq����}����q�rX�]�"c ��^�J��2�����ݟ���O�͛PA,q�:�/$YP����-��|��������2���t�h�N#�Ǐ��b��~���"~6���aq��yx6�n)_���fx'v�ao.\C�k�Ǆ}�tF�W�1'����
3�м�1#���q���3B��*w���k�t�f��T1�"��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$c��X	��MUt��!r�
C���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��N���8@�we ��g庌NA(fۉ���$,��F܂d�ۤ�m�>!����J�Cp�������s�`�|O�\�+�q�� 6x�@�	�x���!��z3�:��c��%2���ʏ!	��c��*;̊���z�1[FQ������-K��s����M�;䌚"\�w��V�)x�?{��J�SqVE�e�H:�I0���ԏ����[���Г�D�i�^�Ax�`Vk���|���sHT�f��H��@!�#-�[ҭ��F6q,/��h�`N���V�I�e!��nH�W�l,ѳ��=c�f������C;��?��QX��WG ��BE�r����`;�nQ�ǡ2�!�7$��q�e<r�4^i�u�J*�Rs�0�|�:���@�����\�H��/Sg� c�Z�qV����Eˎ]":V�C���*DwS9<~�p_�X����)ͶG�q�5�SU*�<�)��z3�:��c��%2���ʏ!����>2{�}����q�rX�]��C`e�n
V~$c��X	��MUt��!v6�RMS���t��B�F�4"��B�*�A���ۖ��<��Ze�C*y=�_�n�To�[>/�®��N���8@�we ��g�n�J+s����$,��F܂d�ۤ�m�>!��˯����9Ǖ��A�\>W�/Z��B���[@���[��QPw��r|��߇(���м	I���������)��H�'J!0��A�6x����V�C���Ul�ٻܔ�ߎ�
1y�A_`OT q��Ko.g()��ikp���H����-��԰�3�I))����A�m�(�A��PmP	�Ȟ�����hLKWਠ9V�-^֬�lPCrM�Zc��qP�U�&�De��2Q�����ݟ���O�͛PA,q���R�*ؕ��A�\>W�/Z���N+~�{-M�O��~�X������<�N������ᴶ;R���F^GQ!�сn����+�Y���� ��@s'R�Rw�)���$G����N�����,eS=�oA��$�J݃����t����9��b>��X����)ͶG�q�5�}�t�ё�F�]	
~ao.\C�k�Eg����0˞����Ti�^�Ax�`Vk���|��܍w�S}��T��̪mMUt��!.���9fj�}�Y�PX�)��s���}H]�˖��1ҙt&H��I����8�����|I]��ם�y��獶���_�(�X�0\[�^"�z�9��IM� I0���ԏ4tv�l�ν�s��U;46��R��O+'�tL�UF�ՁS�Ut�\�|��������2���tԷ���t���3D�� <@��fG�H�*x�߀�q��Nʉ�(Q��;��b�=��|�L�@N|��|(F9%2�8����Ѐ;��i2n_��s�I�A螗�L�͛L�_�n�To�[��Oy�,rw�&�z<a��N� �#{W��:�?"�����JﾥI��ǌ~n`��R�	iT�O����/�k&������&�4z�dט�w������Gl�N~)�jA( ����_�h3��{I��Z��H1c�f���2�خa�>����n8���ٳ��溂�ZI8'��@I��'��q�2�_:��p\I��� ±�sR�{F3�_� ���p� Z���I��'����0i������;�qW�;ۂ��IÙ=�H��M���8 �i��)#bB��G�_��V��6������L~���C�4j�q] ����)_��5�Y�w����K�@��|	0������v��I��RhF��G����FX�,4�?n�=���W�s~��y�.l�8I5�%�l�{�a�I�.��S�[U�JP.D���]�Tk)������7A�SWb��T�Q5�B�Y͘�͉�I����D��õ��Kht-���3Ve�=�k����v��'��Yf�Nd+l�Yҽ֗��)��������Z��e��I��CqZ��v�7
�7��K���I�5����`K��fx'v�ao.\C�k�Ԝ�6NzL͊�q��]� ���_�hbvk~�#xǩ"�4s2nQ�rVwp齰� ͌4s+�ny�T(#�I�I))����A�m�(1#��Z�����XP��ȭb��v݋N�����Yգq����%��/q|��]��0�ȍ�x�>c��w��'o��b9�����)^s{����иܖ����S���0i���R�&H�����̜�I0���ԏ�.fOe	��f�QaK�P�y� "X�<p�Qd����uXӦ��9���I5�4`UV#-�[ҭ���~����'n�^0o��N:�@?u�hk��Y��A�m�(�֟">�#��"5�o٥��e���\$���<3�zE�-~}���%��/q|��M����A�m�(X@�9斻	zL͊�q���Z����p��R�}vJ^ �5�h���.��&GZ>.�0S'� �ު���g8��� ӫ/��m�a��ya�X�Aj����U)+N���Ix���Ka�R8�ܻ��\�vś��Z1`�N�ǁ�f�T�B����$Ů���zւ���MȜ,��Sq'��kA&4,� ���3�ҺIÙ=�H�8�>r&���R�}vJ^�k��76�Z�u2ۅc�t\�<��C娤l����pQ/7j�F��2JHn��z�C����f�SG㴊�?����q5�n��۷I��L}JB�1:���0_hW�D$2���7 E�B��uѯ�O�x z�Jm]A�/���s��m�z����9C��,ў1�ˏ�~ǹ�z��hbvk~�#x��%��#��#���F��-��j��͌4s+�ny���.�R4������˫p}�񥒐&d�X0��A( ����_�s꘤�I��-�3��&Oa9Y֪{���ɖ?��_T���a�aq�������9X�.ᬵy��j��G#���%��/q|z��V&m�����'�>z�/^;؊��yɁ�U�4];ˍH�N"�l�V�����1�so��d�a�e�����c��%$Z'RpW��eB�1VV�zcj[�?�4��ic�v�QZ�?��
���O��5�ϟvзq8�Ј؅��FJ��v%a��!)�����f�ƳaBA�u����`�1�aw����̬��z<����]��#�z2�ŕ�+��/؞�{��^:���KH��˂�%(@/^;؊���)pL��1x�]�V����ߞ�K� �0��k{.Dt�0�Fc�<5�s z�����˫p}�񥒐V�zcj[�h�]h�V�jsUD������]��#�+�9R�зq8�Ј؅��FJ��v%a��!)�����f�ƳaBA�u����`���?ͮ����P�y��3� `A��~E��=��*87���l��P^���֮���"xC��-�T(u	M^�.�/�92JHn��z���7帘��3�=r����0�i/ȇ3
�v�v-}�	mpŴY����;���NA��sm.�9I��'���p�+m*��"Ϩ+`�|��K�z-/����IÙ=�H2�LpOJEl��Q�P�]zm?9ۄ��d1$�Q�<om��7�4����5
iEE�Gg�{�]4�W/S��8(�E���Kt�+Yi=��o�IÙ=�H�R���w(��ES���v�8:��|`��'J�	�LÆ��E� )�&�2���O�}��M�+�'�̗�����L6)�Ey������i�s̍�(��g�{�]4�W/S��8(�E���Kt�4O���x�1��&vl�JHn��z��p�Sg�3�z��SR:g()��ikp���H����Q#�?���;���N%�:+W���݇4�a�Ȃ�u�.�1�a-���7a
��r����~v���b9���eSܥOH�&q^�`
�c��><�$�;m#%�S���RY��.ZVRѿUJ��\���^�W+`�x�oP��@t�&�e�5
�`#_G����q�41&q^�`
�c��><�$��;mQ��8���/�>�W�Y��G��x�&+8@V����L��\�E�V�6IWJE�r���秹�3I^�v�%j����L�de��-@��F~*7���&�_���/���l���F�8���/����RY��k�:A�	S�r��AR1<�N�؆�B��W+`�x�o���{��&�e�5
��Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX�����/��&����H���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8����ٺ?�R�^Ƒ����"X��[7��Eb�qz�^vh;:��B�5{��
��D&e�2l��4�y��ɦ�k�:A�	S�r��AR1<I�0�f�#�Օ��qvdЧ^{�j�g��U-�e��`�?��L��l�%���V���3{��m��rr��AR1<�N�؆�B��W+`�x�oP��@t��4�u>ο��D��$t�գpP�l�L��M�,���	N^�U��ߋ��@�$��Xo��GR��)~s�����j�|��IÙ=�Hw¹��<d�7�
XǺ��g�,P�n!K��tf��
_�n�@/%{�;���;�L���9�D_�3���U_�+X���=ў@'���Xw�j�7��ct�:��RE�QS����>��"X��[9R�A�m���(������{�VwtZ�+�������I?�"Ƈ5����`Ke,fi�U�ž�'�t_�GZEh5���'n�^0o�hŁw:����v�8:��|`��'J�	�LÆ�c�9ʼ��$�G�nJ `1	�<�����!�F<�+P���I��ž�'�t_�B�uʡ p�m~|��;~7����WF�r�f�t+Yi=��o�IÙ=�H��w�K��b�����(`��ү/�O'�=�eX�
\;�M +�gf���a\Y���c_����+#��.X���*"v%)��Qcm hP"G�wk�P#7!smWF�r�f�t���ӯIJ ��`y���Ӻ��C
�y�yi
Y�2}�<��b;�B�W@:`D�h�#�*"v%)��2������1��5�;-;*�7��\@�iz��nVub]߹jGy�ˆn��?g��s>�=�+\{Yh��|����=%+]Bo�A;h�F��O�i��Ե�"xC��:��]<}J���K;�{�&��Y=�ĵ�"xC��}Vq$GѲۯzD[�'n�^0o**�ХM
�?�p�5��9&q^�`
�c��><�$\@�iz��nVub]߹jGy�ˆn��'5 �{B6$��O�&��;�L���9�D_�3���U_�+X��?<�����z��d>3EKrM3�V��g
*C�c�.[K��m w�wAk�Ya�����&��Y=�ĵ�"xC��-�T(u	M^yM��5a�)��\�v�g�W�I�H�¦ʹ
�֕v�՗ɕ�a\Y����+���LQ�X�E��uky�ѱ.��tGy�ˆn����N��+�j|j6� �T˳͠m�xW��-#��klJ�V�Gy�ˆn����N��+����]��/��=6�s���"[��g�7���ìT�T�D��ao.\C�kWUk/y@)�'n�^0o**�ХM
����@tD ӫ/��mR�MP��G��E�hxǉ �Ş(�/�K^b�Mc��_�j��i}q�^r�m�����ч��Z�Bh��vJ*�Rs�08�b(��[Nێ>�d�|Z�j��?�N�@E�Vm�.����O�<om��*)�)q	�cY�~�"���ʷ�J�	�LÆ���#��5q�ЀY@ɓ�M����*��1�G�p�Pv�?Rr�f���,(���B���̴_��EI?�R��n��am�Za(􆿳��1�Q�/L�9d������K)zum��3A�)Oqy�&�CA�o�R�GI$��ǂcY�~�s<��MR�vH9��!e�<�:ӫ���m����������p�m~|��8yL2�����ތ�1��\�vŶ�T���Ĉ��r�]@s��I�λT�v��1���2���I��'�f�Nd+l��_]���T��\�vś��Z1`�x�y�Zglё�H�a)ߤ/؞�{��U\��,�v��|O�\�+�q�� 6x�@1#��Z�����XP���f�Nd+l5����F���
�v�fp�m~|�֚?��]t���Ʊ�_�eD�I�1#��Z�����XP���#���1���Q��ǺΕ�|7J���U�
wl�G[@���j|Z�a�P�Fpwe�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cUL숬W@P͊Y�7#�xI��;mQ��8���/���>k��HB8�	Sc׿Z��A�.ݵ��]}�����ǩJ�9~0X�,4�?n˩�Ϊ����+p[a��*��O�t�L\ ү���f�qNS3�I��'���?"3�m�����h�n*��(�1#��Z�����XP���SG㴊�?����q5�n����a�-�I))����A�m�(Qce��ȢF:����Į��KH ���"���e�S&|���BY��l��=5;N�����O�%��/q|O{��%R�A|�stUy��DbY}n��^[_�e��IÙ=�H��=!ߎ�΂l��=5;$]��Af��s �%��<��x�>c��w��'o�c�.�09m�����
��\�H��/Sg�w��'o�V���"�V���Q�9eY��b��(�F��`JHn��z�V~�#d�	���}�pIɽ�Jz_���0�m��Ϥ/؞�{��ޝ
������U��R�~1#��Z�����XP���K�|q��=H��6�����рӚx��~ ������D>QJ A/��g�đ\e�y��3g��y����Z�� P��\�v��\aьIR=A�;�֋`NǙ#Y\��?�l~�U�{}��*���M!󂋷�(����C4'n��=?���͞��>(�J5l�����+���Zz*��5����`K���}0x��F�ԟ���Gy?�p����=R%�Kw	�F[>�y��W�}�|3����"��q�p�m~|����U0����d5�:�w�+���LQ��U�"����92<ZW`���<d���;����������r��E1�;�>�t$nXZh��\���'����%�a����ǕGF��a�1�Z���=�Ln��S�W�7����KPy]/�qF��G��Q���'��{ �=�%�*�]�1ꘐ�݇4�ae_�d
���ݪ��1#��Z�����XP��ȗd�uY��K��T��p��`�Q;?�͆�%l9�e\EV	����w1�'l�%��>/Q١Ӿ�$d��I��f�:*��v��o̙HxҀ9�@3��}th��.)rL!��di+9DjuU����Uxc���ł\�ԫAJ�T�q?�R��nścp�B��ҍ���������zP�����1#��Z�����XP������0/�e��9�S��8�U]k�(���B����_T���a�aq���U�n;p�m~|�֙X�D��U9����u�I���'����=���a���œ�,���%�a��Ϊ/�^�`0M�/�s���'n�^0o߲�}�{�%��/q|;��c���X�����w�JHn��z��S3W�K@8`+*��A��}Å�S�9o��*�w�+���LQ��J'�!�����qԏV���"�V(�b�|�5�ȧ��i�}��ڻ1�O���-�SIÙ=�H&I�3�b�}�IUr��Ӈih�|���he��G��֥��ع��&j	Z��pDY~��G��5�j�B���� ����H�ʱˡ����V�Ů���z�X�D��g�S�<�c�V�f�;���'n�^0or�.@,j#-�����1�����.��4�F1����������kר�'"I������Q�2i��e�����H����8�N����<�js��0<�%��/q|�-�(���$3 ����.`�$�4zL͊�q����1�9�\I%ji�7��
#>:��� �rmd�&l�����H���sJ*�Rs�08�b(���os0c��ZLN�	��2�V�a��h �x�����p����wя�JHn��z���7帘�f,�s��Zrt�\0�{�ms�A���S\�H��/Sg�w��'o����v�]�Uʚ7�ܩ�.fOe	��|�T������~RK܃��hbvk~�#xeayA���r�&U������G|M��'N�KR���c&;g���!a�`:O���1#��Z�����XP���B�m�/gV�gK����1�*S�b��v݋N������oV��'wNF:����Į��KH ��*PX�KL7��Ѹ��R["��J*�Rs�08�b(���zY�l��R�}vJ^�?�1�{{L	�0t�VW�ȏ�k��a�s+�ҟ�r/�^��D途�؎���ɿJ�:9�2����rR#K�pl� �PP��ƿ�c �B�dH�7DR�i�Ρ��˧T������X�p0�&�����Q�a5���nXZjwi�U���Mչ�����Y��n�Z(Ρ����u�PBxN��X*d��Uf�Y9��_QzMy㥁�hK�'�njVfV)~�`V%'�\�*�c�-@�dƟ�&7��"=��Nc�&�Ia�΁�a�n��!�`�(i3�n`5�fK��@5���<ZJ�hEc�>���gZsT)!�`�(i3!�`�(i3�n`5�fK��0z�cUL(���r�<Uee�N��������=��*h}Nw����
�t�J8I,t�A9�AD�of�7���A3�(N��㎏qló��@d�������e!M^С$���v�|[��5�e`��9�����_�t�y�p[���d�٣���������ݹ�0�����7=����2PW�uD}%V�����F˯�+)�F�������T�\ ��i3�|)sՀ�23
������?�`d�ƇBHx\�'���Xw s4S�'�i��`�z��Y��)�?Z�����1�����NR�^Ƒ����"X��[��Q[R�75�e`��9��əS\��O�=�Q���d�٣���������ݹ�0���f�Nd+l�Yҽ֗�?��}�ͭ��I7��-5��6��	���`y���pzl��a�a���k�_�aY��|�p�6��Hh�]�!��M8���	D%��_�ͅ��I4��欱���j����B�:|l���������CyW�f�tR�wX��J�W��7/�2��2,��g�ܧ*y�E����F!K��tf��
_�n�@/%{�;����f�kN�ı��U��+�Xa�H(�˕-+��B�G����n9�}������ݼ��s�G�7s�9���on�-�6��
�jW��D���M���o�G�m�?%^�����I7��-5r�p =(�a(􆿳�ټ*w2�56ݓ��E���vj��$L�>��07s�9���on�-�6��
�jW��D���M���o�G�m�?�{|*�"�Vx�%L��W��_�ړ8���/����,DTc�~y��i���n���gW���D��g����H���	N^�U{xN��i>r�<Uee���R�}vJ^�k��76�a'�<� \�� |+vܽ�Ϝ��*@&���+�J��Y�{'%s���'���ը��_�\G��4�	B45ƃ
ᾆ�x�T�\ ���|.�Tӏ�푧)��������Ē�LwʅK�'���Xw�j�7�����0/�e��9�S'6���;8=�g��U-�ez�r�6�<n��nN�6�ϟ��n`5�fK��0z�cUL�8� �,�����°������R�wX��}�
�?�r��gGr�`@��q�'���Xw���,D�Z5���l��Vm]�]�!��8�$LQ����ɷ���/s�1��p"�,�>E��P"G�wk�١��	;q�J�� m�h�5,Wlr�r%)cA�z���a�R�wX����K�Q�4br��yO{��`�
q��T�ٮ|�,
������|�FIsŭf�ҿG�p�PR��{�&�8���/�a'�<� \f���ѩj�Q%I4���kN�����~\[$Q��
�`�ю龤9>(�vgH����8�Ј�&��g3�g��U-�e,%�0g��Յ�HN9�VTҝD!u�E����FAԢ�a\��F�dH�Dj���G�Օ��qvdЧ^{�j����#oM������ݓ��E�S���%��ì�u"4�E��b8�"e�<�:�t8:���M#�&���Z02t��S�D�����X���*"��Z�w�l#���i�ɷ���w�kkr��$X� .�/��`~�ߪ ��e��R��!kr�]Q�I����y�搲)���$:N�8.����6�Y�r�7"�p+�@���5���u�L�xZ��j�
�iB{�Z�_�+��tI�F�;���Nk��}�y:�8���/�a'�<� \�;�m�PV|1�#��d_hs�^Ξ�N�@E�Vm�.����O�<om����`��Cg�j*8a�.&�}�z73���߈�90�z��d>"I�`�c{�.ᬵy����5�t�׭��K�Q��萬�]Yݼ��4cGy�ˆn����2�-���J*�Rs�0�5�N�~u=�����z�Hi�����J���e͉�Xk�b��v݋N�����5}	��D&�}�
�?�����}�)r����'���Xw�j�7��ct�:��RE��W��_�ړ8���/����,D�=P��[��1�U���]�!��	Ǹ�y85��L�@��f����k��$A�h��+Fen����9��0|~�LL�a(􆿳���2����.\�#$�ÙA�B�r���n`5�fK�\w��0]7��"=����B*�9u6�|�fF�AԢ�a\�y�T�g}�Ӄ�Q[R�75�e`��9G$�ء���Q]� _ό���.�}�
�?�ʬw�S��зq8�Ј'���Xw���,DH�v�����] 1�0µ�]�!����w�Հ�*��9W��}�bo{W7s�9���o>��l%i�-ݓ��E���p��b����b�g�Z鎬�������(���8'qG%��Y�7#�xI��W��_�ړ8���/���T�/ʍ��)�`E5Xy+�Mk!P����!�`�(i3xZ��j�
����d�R�wX���7�b���������j𛚆z�Ji��U,�(�)8���0y�	�z��SR:g()��ikp���H���F`���G���`y��������5O�KlAP}k�`�B7d��U,�(�)8�}�Y�ןw�8���/�<F� ���Ձ��H��?��m��M�h{;��Tb���/؞�{��No�JH]���oAB�E����F}�=Ll�����&}0�@V���"�Vh�j _ש���yb5���[b�I���Ψ��F�wc�}�![B�
���}h�[�u O	KA��߇5����`K���ػ�T�p~z�r,J����!_�IÙ=�H�8��6�O���it	�Tߦ^Cg��)1�q�ܲ�xΠ��yGb�dW���bhbvk~�#xnůc��o@h�5,Wlr�r%)cA�-��h�m ӫ/��m��?�4D+w�����������f�l��=5;���wGu�ܝ�s2����˨(�V�֪��o�� �}��2m���l������L��@X�hD��$_s����z2�v�~�g��27�*Y=���į�4 _;��i�1@�f=H5H�n��cM�r�z�IF�˞�Bxη�H��:�-).^QQe���b�q��T�ٮ|�,
���h���J	�0�ȷS�J����Xa(􆿳����d/h�5�G�GY�)�}��EXs70��lJ��튝�b�Bϱ���w�K�	�<���BSG�p�P��<jV���\�H��/Sg�w��'o�6��T���7�8���/��Y�r�7"����#!f��$��
�5L��m}I� �-5$�sD$��y�,��1��'�al��p��g��k��i�l����@����gG1N����F�m�^�r�Ϊ�?��(��I@1���t$I+��f�kN�ı*�7`����M�Z���	4����/����DP֞ �X�m��{�Kd#���x;*�}Ւ�~ܔp�l
d��U�9�r�<Uee�N��������=��*pzl��a�)�O�=�}���N|�H�eA ��	�.l�L��M�,���	N^�U�}�g7�}�ξ���I��RhF���9���x��a'�<� \��y��`��0Exz҈��E�5��
��D&e�2l��4(�de�QV踫g(�r�N�ǁ�f�T��p_U
#W���g
����DzL㡉�&�@�}7�q��J��v1a{J��Ǻ CN��a\Y������ԻV8�I��RhF��j���W����T�\ ���|.�Tӏ~�L���vi��N�Na����g�,0 �����r�&Ɓ>i[�ͧ�?Y�Q��ǺΕ�A�m�(�hU_��_��`y���pzl��a�	�_��:�����C��֑xGV�^ɡ|z3�{.ZVRѿUJJ��.U��۩I4��欱���j����L;Л��������
�CӞD��gn�=4�D-'��7�q����d�`��	Q��[�$��X�H
$������Y��)�k������a(􆿳���Qs��������DzL�-��;���iA'R�	���i�(r]m��p�ռ�[�$��X�՚��l��H�/�n>�.-,��Sq'��_�H����K�Q� ׻�1��k]m�����9��|����⾘���c�SD釛-���>T�=�	o #���}�pIɽ�Jz_��|.�Tӏ���\42U|u='�c�-��;���֤���n�V ��a�'���Xw�j�7������7���{r���x�] %� /s��EB�w���%���ց���=�g��U-�e5��e6²]�N��&�#�(�>^�l�'s{	�h�v1a{J��Y��V�AԢ�a\�D�����R�`�|��K�z�
��vK���p�+m*��"Ϩ+`�|��K�z�Q��Y����Qs��������DzL�C��(3���-��w��k]m��F��w�6$�Gy�ˆn����N��+���o�u��"����DzL�C��(3��7�q��J��v1a{J�֋��DO��'���Xw�j�7������7���{r���x�] %� /s��EB�w���%���ց���=�g��U-�e5��e6²]�N��&�#�(�>^�l��e�eV�F��zF�ۗ���4@{A�L�de��-@��F~*7���&�__y�� ��j �0tw�*AI���J�V�	l��T�\ ���|.�Tӏ���\42U|u='�c�a����gW��_K��� X���/�K^b��6&��^�<��J���_]�N��&���3�L����e�eV�M�z$��P�;�G'Ǔ���"xC��}Vq$GѲ��W��mTS{lGD�V�B���q5�n-�@�4ڧ��~��r�pzl��a�	�_��:�����C��֑xGV�eU���("�,�+rr�N�@E�V����P3���2��:�kŔ=�	o #���}�pIɽ�Jz_��|.�Tӏ~�L���vi��N�Na����g�6���Q,|p��<_^H�z��d>3EKrM3�Vy�oY�E@���Rpy2:�׹��t��`�J9�S��˰v���K�Q�3R�e��ł)w���m�±��m|J�}�֖�gH.��2}�<��bl���>s�q?H^��2y�搲)���$:N�8.����6��J���_�Oi9L�:�k]m��,�۞��	���/y��g�'b�t	�U���C��O]r�<Uee���R�}vJ^����`a��R<�����á�~O��L;Л��|#9���b!��u��Ɔ �����Vd��[�l\�`�|��K�z��@d��ץr�&U������G|M���t�2���*!��kѶ���� ㏞ �ب*6��X#���=0Q�9oÖ�"Hi$|��ڵ�)���ͦ��^`��dg�M�q�9�}P�uB�b�#t����n>�YR��j�DI߃��K�+���w���QȘ�d�o/�d��7���ìJ���m����g/��`��ٞ�R̕q���id I�pzl��a�N��	�Ȓ�cЉ�MOc�����2}�<��b;�B�W@(��T�[�=�5x��j|�>�OU��9��]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e5��e6²�T:���V�����,Ǣ� ��^�:Z鎬�������(���`$�P.eE���lC��U�T�\ ���|.�TӏU�m#j[W, +$IA ͒�ښ�l�L��M�,���	N^�U{xN��i>�/�n>�.-,��Sq'��_�H����K�QR�Xe�������(2���􇃬Tk��A3�(N��㎏qló2u?r���Y�G�˱�ߓC娤l���Mq&���[�=�5x��M��%LS�8o�f���k�:A�	S�r��AR1<]Q�I����y�搲)���$:N�8.����6a'�<� \|���yB�+�kv޶Gl��C*�󅒣$���:�kw�j��,�0�@vV��
��D&e�2l��4��a��se�`��ٞ�R̕q���id I�|��{>��e�t�b���6U(�<"s����&=�rs�i��O3JT�!I�T�\ ���|.�Tӏe�t�b���6U(�<"�%�2C��rs�i��O3JT�!I�T�\ ���|.�Tӏ ���v�l.�
��ڋ��Q]� _�rs�i�CЎ�����Ɛg)x�D�����X��Q��Y����Qs������T�e�V0�� ��vзq8�Ј'���Xw�j�7��	3i�\��׹��t�M��|S�/����Øf��K�Q��`�����!�`�(i3�d�٣�����6>��JX-�ܶ�0����K�� ��^�:Z鎬����Y�V��#qX�9y��"Y����8eZ鎬�������(���SG㴊�?����q5�n�@qQ�ܩ�8���/�a'�<� \纅<S�O؏����:aޗ�U$�'���Xw�j�7��	3i�\��׹��t�M��|S�/������������bpO؏����:.Ɓ�dd?QZ鎬����Y�V��#qe�t�b����t]������ī��]�!���1����mA<�}	��G��[�f�]n�"��V��d�٣��c�A�L'J����l�!��G��+�c#K�e m8�8���/�a'�<� \<F��̎ÆLx�A�B�m@�:\*�Z鎬�������(������aU�����w��T�\ ���|.�Tӏ�'�ŀP��3B�\G��ﱴ=�]�!��	Ǹ�y85��5m*�Y��g�S�<�c�!���X��`y���pzl��a�D���ƨ��u��u���� ��)p'���Xwa'�<� \f���5���w_������8T��]�!��i��&�J@{L�'x�$vcH���K�Q��2�����z��I/r���+b�a�&!9�q5 ̬����b9����Z[Zz�! HڜԎ���J@{L�'x�$vcH���2�1L+�&!9�q5 ̬���M�8��;[�(��Jx��'�!�Ѣ$X�jl�N� �$]2�/.ePN6����(�;UW���g��'�|v*�n�6��.���I��N�\Ӽ�gy�A=D�!v�w�u��.tƙ��3Ve�;�0�XǷ
�J8����d��MT�D�9�.g^�F���p>�����;mG�����k�}�m
ˈ��$����q���w*��	�a��������t��P�mjS�z�9U�s�Z{�=����X��-��sޛԪpP���4�?CZ=x 
~�F�踫g(�r�N�ǁ�f�T��p_U
#;��|B��>>0j��Ih�	�;��J�����M���R��ӟ-�F���ˏ��Z��zf	�$NT�I���I���C1zh=E�g�N�������S�_
�u��Yx�I���I���C1zh�6���Q,|�rHYSڣ��ǡ�C�a\Y����+���LQ�s�xV��8���&�@�}7�q��J��v1a{J�?��кDO�,\���ӟ�X���&�@�}7�q��J��v1a{J�d�	@f�u �U�N;k��!a�tc�&ck���>#qBK"6j�"Hs���ٚj�ώ ���]q��J��56�f�s�G��J�����M���R��ӟ-���4�&����Z��zf	�$NT�I���I���C1zh=E�g�N�8�dEm7�w�kkr�I�;(�\��8p���uAԢ�a\�DW��E��q�����C��֑xGV�eU���(�CK{D�sss2����`�|��K�z˦9��iժG�p�P���ً ��3R�e��Ӵ�"�6j��;٬sf.�5^����r���zk2�����n�۴�.�<Mm1���P�|T����E�E��3�L����e�eV�M�z$��P�Ġy�����l�p�H1�a-���7a
��r�$Dc~4�A)�V��/�c����sL]~цt�U(i��[���P��d��MT����k!Tޙ�ǗL��	��q�©�����<�������~s���^��{�)�V���x�l��1:�N�*�xA�sxW�O�Ji�];���ss2����`�|��K�z��u��n�����\{F˯�+)Ƌ��_��F˯�+)ƾIwL_̫"���	��,�nY[��o���a5��EfVNN{s�ܱ?'ÔhNVBN���
���O��5�ϟv%[�1�wG�}M,�d��T��ޔhNVBN��
�5K�ƠX�L-�.n��B*T�gR� �ұ�X;p`�gR� �ұݼ\suLﭨ "5�]�$�`V1���n�|����Y�{'%s���F���gn�=4�D-'��7�q������X����}��uJ�'B�ɏ��]�!��	Ǹ�y85�0+ע 5N�I���I�����O!ݨ���0[4���$�d����==�h�f��z�taS���	h	�/�����	p)�O�=�}���N|�H�e5N�	�k��@����:_���oC�����8y����
f8�|s��_F�k-�H��b��:��6��<�]�Ե����)%+�O�W,�P 3#4���-�� ���JH����8��#I�ND�s���H�V��^�5G�����&�@�}�-��w��k]m����8��G��,\���ӟ�X���&�@�}�-��w��k]m��+qO1U�)�#qp���W/S��8(�E���Kt�n ~���7��3R�e��Ӵ�"�6j��;٬sf.��ǞZ߻��^E4+у��b�Bϱ��3R�e��Ӵ�"�6j��;٬sf.�r� F�3N����Od-@��F~*7���&�_$� %7䨁c����t& ��i�߬�F�<H�n��TD��-���G$�3#4���-�� ���JH����8����F)�~����H�V��^�5G�����&�@�}�-��w��k]m����8��G��YN
��)es��S���.�<Mm1���P�|T����E�E��3�L���'s{	�h�v1a{J��>�_��� �U�N;k��!a�tc�&ck��Nx�P��A���TaZ/����>��i��N�Na����g���\v2:R�S�yN4�S���%��N[�[^��k����x�xG���۵z ��gn�=4�4�	���WdM4@��&����˶p�0u�xs�&q^�`
�c��><�$("�P��_��3�.�J�|�+��?�d���&��$ͯ����mѷ���V�象�;��_�=�������+��T����oGo�Z�������/�)��ɖ`ۺ������Xc�F�������ϲ�>e��>��0��E|�,VK�5��&q^�`
�c��><�$���E������Kp&�w�%b��G�w�Iſ�Κes��O�h�S{�5��lW0�c4�j
Թ��~��q����U����*]S����l��))^{?	�c;@D�
��Io�p��76,�/^;؊��G��𤰇X]��U�I&�j1b�jT�.���I�]�Bb���{��¸�m�B��d���m l�o�@`�~�&E4@Q�/�9��?xsl��)��'���Xw�j�7���3R�e��ł)w���m�±��m|8�����F��A�����~W��� �A�J�e�!�c�A�L'ӸT�?��i��N�Na����g���\v2:R;�/B��[b�0<��U�%
�bql�d_b�~�`�S��P����{�j%a}�C}��0Ex�3,����W��2�H=�m<����6U(�<"�͊�������?�Tl���FѱTW%#3?���*��+kt�Oz�Pa�(d�b�W)��/80����)��K�Ԟ-zq��Qo����Ԟ-zq�r��iN�!���5�Nnb�k��g�\k%��N���,Rbc�z�F��Z��/�+S6���N�@K��SRt�1q����C?�+H�~���g2��\�b���]�M�v b��0�s������mroL�J!�Pip<ɯ�n��\�XH�@Pψo���Xgn�4�K�&�|\��t��Hg$V�����EyV�Ӆ7���L�УΛ
V+��W�p��)8"O�,��_u�wl/���(���eC����9��Qm.�̸��Kv�BB$�W%�)�h`��{E�T�`>��6�����#c�%���>M�-��<;:��t� �?�w-���&Y��V��'&�s��M�Ǫ��P`$��*�!��;�B�~�{�Jt+��F�6�B���Li�����E��u�H�h���^��%�fE�DĒ^����' ��Y!�Y;e�iK ����)c�g�0�u�'ž1�|e�Ɵ�s�܇��9�R연e�E�k�\D!��,b���e��0�U+�qbp@��\�G����11�����c�����hX��WG ��ASU�
T_�mS8<�n�5Zbz�Z��e�E�k�\D!����_g�$�����[m��3R�e�����v��a�Ż�&ǥ��a���F�LFC7�5$�)�vx8�t��_�t�C�k"LB������ׁFy��_y� '�u�12�'�{����Md�sω��=��m-���T�}ɻY~�y�����[�T���Ӫ!��˼�v��j��@	�<��k]m�����9��|0�rI+�ܡD�:F}���V6��Q��&i��N�N-��;��M�z$��P�^�6�V���l�p�H1�a-���7a
��r��s�]�x1~�D�#�iA'R�	���i�(r]��0�|�ʮ��º�>:��_
�u��Yx�I���I�����OeU���(x"��!!���l�p�H1�a-���7a
��r�S�B+����;��|B"�2�,.�Rg��L�*�ZRk�j�fXt�U(i��$�d'X7���2�"�G�p�P�(��Iw?�d���&�B��QY_��֑xGV�F�m���}'!��/����'���_�����o���F��!���Dڋ��mhcA��짦���O�ʦ
���c�v�_����J�����&����˶p�0u�xs�&q^�`
�c��><�$("�P��_��3�.�J�s�xV��8a����g{A�dha#4��������o�^Һ�i�<�~�yا��=tu�Iy��F� ��N.i�AԢ�a\�DW��E��q��u���'b�'=�(J�}�֖�hKBi����1��-+Dk��!a�tc�&ck��Nx�P��A���TaZ/@[�_zβr�j5�{��2��@N�X��!�_Pw�?��?hO���&z��kɡ�ܬUvd���n{�5���6�V(>��uh*�%KJ�	�LÆ�b���[Q�k� �QJ*�Rs�08�b(��,
�u#��!�c��V��������hm���S�Է�Æ�q�©�����<�������~s���^��g��%��,\ަ�Itݡs����0�r<�V��w�%b��Gv����Y���a\Y����+���LQ��xy�'�ӛ�����\����>'��������B�bq��ٙ���O�#t%zY#G)t����G��7������D��t�!z�t�-$�I����Q��K�%�x2f�G)��j)yc�n�.�_�t��*' 1�M�ʦH�K��}M,�d�}}wS�7�}r���՗����ڃ�"��
!�7��?\�����(f����U� �1�}�l����+g�%Y��̗0z�cULj� 1�-��;���iA'R�	���i�(r]��0�|�� L��72�^�9.�JQ�0��"��S8�TkF���㬲���OF�m���}'!��/������ٝ����|�Y�_e2o�R�r��h�f��$;pIGB����������5Zbz�Z�f$n�L��4�g��n%�)eUȯ���3J�~{���Bb�<�kɡ��?}I���]�}�b��~�O&�r�$��3~���s���@gr��r�N��lsσw�kzbp4���o�t����s��G�Ȧj�E��g�Hb~�f��*K�K8����Q�z,;7��"U:@ jG�uh*�%KJ�	�LÆ��5$��?��9|Q�ZyU)x�?{���x.�Knq��$��W*xkx U�_@��D]�V ��Y!�Y;e�iK ����)c���������]��!k����9EX��WG ��k:j%]a6J�ڣ.�����2����b_X�XV�b�z'hۉ)��R����\�G����11�����c�����hX��WG ��������M�h�ˁs����a-6�Da���P�]��w]3k�ul�W�� ,��rQ��i��z����>����:��KY׏�����Mrw�&�z<aSm�6��`߸��S�Ȍ�:Ll~�]��9pq66j�"HsF(��#U>Z���X����9^*5�E&l�z�Ԟ-zq�-8c�i��9�W8�|�wqMYxw��N�u�-���t��P��M��%LS��$E����+�~>�ŧX�m��{�6;���D8��2N!�y{+�4��s��Z���.T�~>7:}nK�c��-k��Q�#*�7`����M�Z���	qb	��G��-������X�m��{��$E�������_g�$�����[m��3R�e����X��9@[�_zβrE��g�Hbz;7��|�G/�V���y"�6���qP�V>tI��RhF��j���W���?�d���&�^�n��Uh��i��z����>�v{��lw	����,Ǣ�����=����,�ǰ���l�{��h�<���@[�_zβr-:S�4����;�B�~�{�Jt+��F�6��Z'� �Y��ݎ-z�;��X�C�HC�|��dq98����H�\�c7����GЀ���A((�����>t�^���\�}R�Xe����s29�2|ev{��lw	����,Ǣ�Пe���;u�4�J��R�Xe����B�%����=;v�g��n%��gn�=4�N�w_1v�V��	��yY�p���G�Ľ����HI�J�@Q�P����ؕ�V��	��yv��r�Y�ԪpP���4��!���缐%�/�<�d�Hk�x7	C���̨�W�Vc�sNL����CQ�f����;zݑ����j�v��3�����5��p�_6d��R@�sŀ��З��:c�<*u�p�Þ�N掤b$�+��mų��n��Uʚ7�ܩ�.fOe	���A���T�T�D��ao.\C�kwFp�����N�"9���b�=�Z{}t�\mc1��^���f�UlM�l�ȷ��>m��Iu�`�o�wqMYxw����S��j|�>�O��Ȧ�R\2@;��ݤ�_?�d���&����C1G�v��X�K�\{
))�H[ɳv��X���&:rJo6������1�R+-h]�pr�}rO�/��^��:I0���ԏ�.fOe	>�~Y�I5�4`UV#-�[ҭ�Pн�cD&�<���#���!=E{J�QF�� ��!�������˞����}CR�Wi���f
hZ�q��a@���-��J�;d�)�݃�(����@�1���Ֆ��}Z�
d~h�7��sBbRt�nr�!m�W�̿�z��lPH�?Y%NtvfI�ihv�X�v�/�Q	m� ϣB�����M��&Y��V��$�r�6��sE���y�q���G��Rs!g�E��V��،���,�M�B�~�)K��a;��]�t3,H9��ܜe��g �q��]����c�o�`R���j>��3�	���%�� 掤b$�+���Nˣ����ġ��,�%X�9��PG"$�m��Y�����|O�\�+�q�� 6x�@�s���s�?�#g�k��R�Xe����ɲ�cz���v{��lw	�c�}�C�ǹւsr⍍N� �J����Ey�mDƝ��0vdLqgF���~v���� n#��Z��w�3�yh�>�#��Q������ssY�KJ�	�LÆ��5$��?����H�V�]cA�x��b�����V�I�e!��nH�W�q3��+���-��Rއ�j|�>�O5X�nd���)�O�=�}���N|�H�e�����W�m�M��%LS�I����5��WS˓C�^�o�3! �����N^�Yإ"i��V��	��yS�L]�z8��8P�j��<�ql�d_b�o�{�R�_�
��[�&�K��A�6�L�t��n�1�+5����w��c��>C��`����|Z!R�߬�F�<�;z�Ni����2�"�G�p�Pڹ��/^�w?�d���&���|��
�|u='�c�a����g_��N�\Y��-#���F}���V6��a[a��|u='�c�a����g��Z]��-@��F~*7���&�__y�� ��j �0tw�*AI����ݴC`�3�<�H��V�[�s���_����J�����hU��!�97��ENҽ��O�ʦ
�[�s���_����J����
i���R|�1�a-���7a
��r�k�Ղ����Y-��V��k�	�"�kϕ=���c����t& ��i�߬�F�<��#����2��@N��;z�Ni����2�"�G�p�P�(��Iw?�d���&���|��
�|u='�c�a����g_��N�\Yfύ-�9-�S���%����g���hZcA��짦���O�ʦ
�[�s���J��sr�l�k]m����ǡ�C�a\Y���[C�W�v/��1h=��]�V/}�j��4�d�cX~|�D́.�.����s�xV��8C��(3���-��w��k]m��oV̲
�r�YN
��)e�
��9��}�����(��b�Bϱ�ɲ�cz���ł)w���m�±��m|�o<4y���W/S��8(�E���Kt�4O���x�'�������p�+m*��"Ϩ+`�|��K�z��l��jV��	��yv�ʯʗ�bu�rd��t�t�#�(�>^�l��e�eV��֤���n�Ҭ�	�
?�Y�{'%s���F�
ɴ��z�4�	���WdM4@Ȏ�U(`�ȕ[n���"'��l����C1zh�@	Ŭޖi&k@C�Ɨ0z�cULj� 1�C��(3���-��w��k]m��v�b��� �7L�a�C�#x����I�?g�f��Qө}�8o�C���7I���ʊR$�ޓea�;y� ,b0V�u�Q��]7K�6�á�~O���-@t�/�W/S��8(�E���Kt�m���i�s���1�R�n� �}DG��^������\{F˯�+)Ƌ��_��F˯�+)ƾIwL_̫"���	��,�nY[��o���a5��EfVNN{s�ܱ?'ÔhNVBN���
���O��5�ϟv%[�1�wG�}M,�d��T��ޔhNVBN��
�5K�ƠX�L-�.n��B*T�gR� �ұ�X;p`�gR� �ұݼ\suL��7's0ۉO�l����+�:��]]t#�(�>^�l�'s{	�h�v1a{J����G�9�'B�ɏ绎��YxP���2�ę�u'b�'=�(9�n���ꢤ�Og�C9r%e�X�m��{��R�k���q�\E��0o@aT�\ө�M��%LS��R�k�����d\��y	��Ƨ�.�u�Q��oY��
�iC>N0Θ�&��GE<Ң�c�����!9�= �m�".5d��ќh~-s/�<�V�QK�}��͢��wqMYxwkDڧ,�R� ,��rQ%����Nx����iV�W�Z�+�~�{9�e��;w��Ĉ���rl���ZJaM�ח�B�Yc��`j��ء�Ch�e���#
�FH!w��z�e�V�{�虀���+j��̅zH�����c�tP����H�!C�Wm��5�4��6�zy�Vނ�L�q$�'�{�ڌ�2W�.��H8���T�=>_5LU�TY��Ĝ(�IyI�Z��7$4 �P����-/��r��g}4����F��ay��E�<VF-x}g���*��g���'e�ɓ�:�a�0'\9�م|Kpn�3��I���s0n3y�Ĉ���rl�n�Ϣ��BW-i+��93G�R�k����Y-)��#�ɀU��S��<�#�A;��|B��a��}��;�gE�w�Gu�������q��X�.fù� ��u��1c��`�D�Ⱥ��qX�����^{��v��@7��z�]M��z,��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ha�Ko��m�\��5/<�KǣDޛ_�.��)n�w�'��Lk}t��]`�L�FZ�1ǿ��^Ý���z4x��x�L�FZ�1�M�ŗ\�'	�?��[Q��Ш�^v��[6"�I�?g�f �H�Z��1]���%��FG�n�t�iZ]XF�hx��G��!�`�(i3n!��i+�ť�n8���L��g�I��RhF��ղ�^=�
t�zg��p��I7��-5l*���T�I7��-5��5Z��·���~X�~���$^!�X;p`�����?�dv��oTN֢&@��&��|��p8=�[Ǵ��p���@Z�_F�k-�H��bf�?ǉ�=�|�)՜�4z�Gb��P�!�`�(i3|w�{P^K���3�<�p�� �&���ç�A!�`�(i3�\�!wn�ř�3�<�p�� �&f��vA<U�=PRpY.[?V��j�cZ)[���F	��7��z_nÑ2h�-]�o�Mt��1���(Gl�q�X癌��� 
~�F�踫g(�r�N�ǁ�f�T��p_U
#;��|B�w,�O�`{�3Vg���j�Txk^�� ���R�^Ƒ����"X��[ow_;O
�xkx U�_@�]t��fg��������B�â2N!�y{+��0Ex��L�.��e��~��������Tg#�o Yt��}��z�S�T�٥��T��?b�t���6����H�5�Y�w���bʺ��)o�N��*M|u�޽�vUM��)�� Ww��Il*~IP���*��N�ǁ�f�T��p_U
#��'8��)���"5�o٥�i��ݟ�^���\�}N�#;��=��ծ�+�� mv{��lw	����,ǢL�E��<U>Hp�y�7Dl�ggi�S��w_��Gb��VH�p�-a�D͢?�d���&�D���ƨ�w]r���nX�i֝�G\ibE�G!@)c�,���M�*��ud�H�A�m�(�����Y���h�ӵeo�;�iD�m;��|B���X/��əS\�R��)�POۭ�نL�t��ni��:$��28��p�!���V��	��y���˳���~�޳^���������G�Ȧj�rZ�0m�\�n�8�Z�Ѽ՗�zϋ�,n�8�Z�Ѽ���9$��H��u�d�ۋI7��-5r�p =(��8�B���ow_;O
�xkx U�_@�]t��f]���^��m���PH�F��׿]=ͅ�J<v�N*�9�c���kb>���pۀ��t�~x����J�u;��|B���0�2u��/n|���<Ӊ��S��A&Qne���J�";��%YM�ξ���I��RhF��j���W���?�d���&��4w�d��˩���.pՁ�=�nlTU�QY�O�5�%]���a(􆿳�k��q��־�E�&�y+�.��.f�Cz瀿3�_Ï_&-T�*�7`����M�Z���	s�����ه4�tZ�=��ծ�+�� m�ݾ-/�;��|Bnf��;�\sf0�s�I�c���;�z�����S��A&Qn�_��1J���t����M~V��	��yޮt
0�_����s�j2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc4�`�(H�Ps�q�6����4�G-rx��� 0v��W5���i7��0!�[�0>�
��`��<�
�d�ξ���Ix���Ka���\�Q�b�#g�k��Ps�q�6�f!��������raǹ}���,*r��`�*Ea;��|B���J����}ָ� ��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϱ�y�Zk��5/��33��*�	�ػ/W��^{Gj��J�1	�<����to��y�[��7%^�W+��W�
cʄѓB�@o��[ea�8���B����g��Tݭ�EB�.���mtPM�^-q�x�l��1:�N�*�x�i�ۑ ��GZ>.�0�<P��C���U��+�Xa�H(�˕�&�C�/�w,�����<v���G�kޮ��n���㬺j;��q,9��n�7�Y����X1Ο<������.��R�}vJ^Z_V�`��n�����������_-�ȩ:T�v��1���e���0߰�%� Zt����$��"��#2ش�T6!�]S>.�ƪ�Qm�(�O��'��+�t2�0�趦���o�Hc�U0�!sH�\`�3J�V����U���@��������=��܄�H#�"8��!�`�(i3;���[���{s�ܱ?'�=|-�e1|E�A�2�1#V���<�dv��oTN֢&@��&���Mڷ�21!t*x�S.!ū�ez��k]m��,�۞��	�rVu,� �{k�h�+|�c�$�t�]�;���VС���u_�P�v	��YY��
�iC>N0Θ��ݚ�Н�bs��2[������	�;�ݚ�Н��Q}mҁ�t����si^��"x?V��.�h%]�lEGV`2B~�={��y�(����1Y�{'%s��	%�Z ���z΃�"�.�u�j��ޓ4�F?P�.!w'L& �N�	��i�(\{ف(�7���<��Y���U��+�Xa�H(�˕��:�EB�Z5�O�%E#PQS��:Z�7G��#{Ձ�=�niF=�xo�n���㬺����D�Ϩg��U-�e a⣃_B7�}�!��N��	�Ȓ�@{2귑�'=��!���wTR}�/�����y���|����'��$zөI��)���W�w��fD�g�9��,Y:�{]%sշ���⪞mf��EYzȧ���2��'B>&�&i�+#c����nS�3�ǻ��d���!iЈH�����2��C�y��1Q(N��vj��$_.��45��U2X��������,�ǰ��������2܌�I(�g�y��6j�"Hs�l��J�&'L& �N��ƟA#F�Z��E��3?�d���&�P��TˇZ+�6�Ƞ�����>�ܫWEFΑǜh����X "
z��_r�e~5�O�%E#P���=J����uS�#̮y�3���;_��8W�w��fD�1�C�#�] �y�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�"��3E9�H�i�e�}�������B�@o��[ea�8���	�~�����F��mF�!؂�����#fr�L�t�iZ]XF�hx��G�����=�-�o&l������g����=�tt"���O�����J��a�U"�^�R@Κ�2e0��Tqmp�AJ�e�$��ݥ�7�����.��4�F1���")d��S7�8�8wGPyn��C!�`�(i3S Ë,�	k|p��z~�I7��-5�B�wj$g�u~xgA�������S3CO��REԔ	�8�����ϲ������i���i�\�>&�&i��&�C�/W����vcy��<
DN��X;p`��d�uY�ؤ��E�����|>U����z~�B�wj$g����d]���GF��a�1�Z���=�,���9^-����m l�o������X;p`�gR� �ұ�BA�IH���O,8(�6k�4d�Lt�2�t4�0 L?�p���@Z�M�g�����X;p`�(������\�LtF�-��{����"q�\E��0�����?M/��k���}������ݼ��s�G�f�?ǉ�=mj�B��V%@��4��]�;���VС���u_�iv�W�O�vA�VG��,m�.٧p$���"��U)���aʍ,wۿ���WG���iZü#{O7��cm�j���X�q�\E��0	ozqP�k��rݾ(����C������Dr�mޅҺ�Q�����*�� �\{ف(�7���<��Y�(��/�h��L���2?�d���&��D�U�2Y�'����2j�Txk^��]��3R������e���%ޘD�P�E6�k��q��־�W+��W��>�:| ǾX�!K9�ҞS�f�
jJrf���QXv�5����%l���V�E�i�m}66j�"Hs��nt)!��(�1�H�,�]� ������x��	A����PqZ�o���ia������v�h�g��U-�e a⣃_B�-���^ncRN�����u_��K��V8��mt�\�l=�L}�[t֕ߝԀ����L}kb>���p����9�d���V��	��yG��Γf�-I�p��g��8�=wF���e�h`�m��6�3٬t�Cc�{A�����M����t���V�~.�
������\���8�'�8")>;h��:.ڥ��r� ���$�Hՙ:Д;�?�́�yuՏ���i����^ʤ�G��������� ����H�ʱˡR�("H��?�d���&�#��`*�Z�u�x�c�lR��~�IX0F�MV�ҁGG�.Mm-;�C>��Ӛ<lȕx��H����Qw�c4~Nr_�mS8<�n�ݚ�Н����*���}���Q�c�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3���*���}���	�g��xE���8����]W&fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��.��vذYC�8����g����<����,�ǰL�[��V���?��;!�G����Ȏx��$�H�ۗ��/?�́�yuՏ���i��}��g�'[�O����� ����H�ʱˡ`����N��?�d���&���腩�z�������:7L����(����C���۵\������,�ǰL�[��V���?��;!�S��9���� iI.s�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�hvb�O*��q�)�`C�G����]'\gWg��	�Z�kfc?�#	*]]�(&�L�xjzӝ���I(͂��-����r�VU���G��5��%�Җ킼nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��yо9�d�L�c]p�5�	$o��Z�_�n�To�[�}�~��l�܍w�S}�H�
+���@�V��lÄ/�,o�9<���F���:��KY�[b%Ɨ��E;Eh	��V�>ȿ��'���#8��c�Z�~p�-a�D͢bP�63Z�tr�VU���G��5���?�1%��?�9ظ��ʱ�_ryhx������a4���܂�`��.��G��[�f�x���w�b��G��58��Տ*=ܑ��y���8���/���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M|]η�� ��������*�:.N{i�tS�SaqZ)�vL��V�>ȿ��'u���MN�G��[�f��!�+n�Zk��tLk��:1j�=�+�T���?�L2��_�#cj1�g���(����5�Z��f��Ո��D��2E�.�b�ySe����1�:�Ω�.�&ʺr����$l-�㰻��V��o5]�Q;�im��ȍry��	w¹��<d���<
DN��$wq����+W���F�^�Y�7#�xI�"dir���r
�a2�r�hr�W�������#��=��kN�*���j�M���rL��GeY�^�R@Κ�2'�̗�����b��Pp��h�5,Wlr�r%)cA��b�'�ſm��'A>� ���.*����Z�j�r
�a2�r�hr�W�:�'&�
no#��٠R�^Ƒ��8!�w� wk���,���9^-���0)]��w�b^X�P�9���TE��a��'�-�1H�3}�?�_�������� "5�]֭�h��Oo��0��7t�%�Z?��<�ry^�h�'f R�X;p`�(������\�LtF�&8�,�#N�)L�*�_�I<�N��KPkqy�{"�i:�gR(]ͅ�y�����5�.?V��j�cB�Y���c
=�2����޴�ik]�f��p�T�q�\E��0</���/�u�[-�c]^�ʎӦ�V�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Y�o��}�����k��h`�H�MPq6.�yܤ�܎~�J���^W�������������_�ft�m-���L%�o5j
�^q�&Ѣ�� ��&6�%�@��n{�\�<:���\���D)�g�%v�=̽�0Բ�ȁ��;�<�h�kIp�#>��QS�����P���LȬ@VYBWh)b�����k-�5����DE�<���5[���������۷�[��7%^�W+��W����#}�Σ��ֳ�m_=uc�cC	�UHtL�#��f���F*�#C(��l�6>8G���n	l��Q;�im��ȍry��	xF���u$J��<
DN��x�8�D"�����ׄ���MK�LWT�/@��R�^Ƒ���X;p`�Q�%�+2����F$f�A�h��+Fen����9��
�{�~S�!�`�(i3+Ώ1;��5�}�]���;�)A��i��G�K$x/��&���&�2�������ȍry��	Y��
�iCTl�������l6���0�&�ͭ�U젩`#�4>?� �1��ɕ�eY�����w6�`:A)*�ݚ�Н���_(x��`ǂ��%D�$��?�')I�wӨj]h����dЕpב�B�^�Mi~_�T����,�ǰ�~as>}{�j׻0
��0i��V���m� D�@G��l��3\门:<#�'	�?��[�%�~�ѢurL�����'G�+R���o��_�Rv�䩲$��GQЌJ
�յ[+8����"sS<�0�zG�������&G�wӨj]h�jsrCm�kE�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l���{$�������LQ�/8n
V~$�(+Q���G�:���f����\�v#i����F/G��Hb� h�ҩ�?V��j�c3R�d�ܦ)�vL�����]W&fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vxI��S�ud��E�9K��;_��8W�w��fD|]η������]�]�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�!I�~��a�.�)[l�P׋��W��+���LQ�M/^���iq�VD�Lg�։�^�c�ؒ)��U��֜��3?�d���&���������oŵE=�k���:+$n�U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�{k�h�+E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l���{$����^V���!ֿ*Y��b"���LQ�/81tSjv�����l��������t�|ݔ�3�5�}�]���&�G"f�x��re�{�W!�`�(i3{k�h�+v{��lw	Sr@�4g]�1�Z���=�"j���b7|#9���!�`�(i3���F��O��ݚ�Н���4�*BqC��~�;ϔW�@Q�kj� *�h,|1���-����!�`�(i3�}������xv�3���Q�j�V4ʐ�}	�[���&�Ł��2a� <4l���dNu��D%0�!�����tg?�� W�hSr@�4g]�1�Z���=��������Z��q�!�`�(i3�������l-�J4p'�>��Q�j�V4ʐ�}	�[���&�Ł��2a� <4l���dNu��D%0�!GmϨ/��� W�hSr@�4g]�1�Z���=�������"xT��z�H�RtV�^!�`�(i3e�v��ҵl+��%�k<.�B�0���;�¬pX��g��U-�e�,���6+�!�`�(i31���~!�`�(i3yo���_$��4,�Q��+�uB;y�F��P��G��Hb� h�ҩ�!�`�(i3{k�h�+&k@C�Ɨ0z�cULE��K3�jާS��m��X�����j�5�%]���=���B�u���P�7� �:5A��p!�`�(i3��jVѭ@!�`�(i3�2��}��cI�*(�'���Xw�j�7��Z�qҪc��g4}���1�Z���=�,0�A��U����z~)���	6�!�`�(i3fĉ>99��A0ok��!�`�(i3���F��O��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6�8���SY�N�o��C�0�b�<�'V��	��y����X�M���������+��QJ�wk����\����|ݔ�3�(n�'�}x?<��U��֜��3?�d���&���������oŵE=��6E_�� �o��_�Rv�䩲$��GQЌJ
�յ[+8����"sS<�0�zG�������&G�wӨj]h�(%����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩ�-��)'�E��ȷ��#o�]�ʄǾH/�d��_�mS8<�n�ݚ�Н�{k�h�+&k@C�Ɨ0z�cUL$8&�{�Nώ�;�|Mg�gqc�e�K���<�ݪ�򈟲�Z��*����%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}Ĳ�y��iE��+�Z4k;/B��.ض6j�"HsЈ0�IMY�����]�]�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hZ��}	�������E���	�������EX��(��n؇�k�.#���2�"�N������A���x�BÛ=����]�Z@i�~���2�"�N�����Ւ-/�;j;��|B@��Ù��Ŋ+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}����F1��Z��Ջ`,9�H�W��`�z��Y��)�gP����,�����J��:���鳖;nSH���k]m�����y{�!�`�(i3!�`�(i3����;q���D)��Y_sĝ��賖;nSH���k]m����{"gY*�7`����M�Z���	����}�ϛ��D)��Y_sĝ���w�R���y�s�7�OTџ�	 >{�P.��L^bV��	��yGn���B ���:t�!��N&��H8�d�~��@*�7`����M�Z���	��]�&�Mc�X�G[����t�T��?E-h��`f���s8����z�:Fa�7���W"�P�K&�c���L��������r$ɓǃl[�Ƶ�1tSjv�O��(���*�̟�1dN�<@Iv��nt=:�֕ߝԀ��`6X���dc�@c�����h��-����;�E����=�O�-v�*_�mS8<�n�ݚ�Н��Y.�~�|����aGl�97��EN�y�JB���PY~�y����o)�T*�c�Q��Ne<��t��y���'j��ݚ�Н��po守�u닓.�`�3+,w	�Af̓@?5�3�Z[���A���ۖ��S�<Ԣ��=aS�H��ݚ�Н��� л����M���X
�g����*�S5 ��ݚ�Н��I��Yq���k$ ���y��lDe7g#�qa�E�Rq���my$�N��o�/���;!�`�(i3烉s)�v�bP�63Z�t��\ Nh�;�P�t�5�� л��5ߧE4�흔\ Nh�;�P�t�5烉s)�v��IX0F�M���M���X��*��� �%����yq����lsφ��<�6�@a� ��fFMqlgʃK�,��`U��B��-ն'�U;|�u}D���L��������r$ɓǃl[�Ƶ�1tSjv�O��(���*�֦�n��{_8�Y��=�}�Vݨ�,bxqX�*qA����6\�4�@�� �-j�1tSjv��po守�u�,l����M?��y�!�`�(i3[�񵻕���M��2"���&�^��v�8:?�'��ᦾ�;���8���U�._�nQ�rV��q�t7�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2E��6x�Hr�6w��]W�I))����A�m�(��ʢ
w�YN
��)e�W�J��H����8�O�5���1tSjv����y��lD%����yq�>f5�� b�z'hۉ)��d�7�q�<�6�Q=��jVѭ@!�`�(i3�Y�
 �vc�jj&��G�9m6�XƤ5_���"~6���aq��k�7� r��L�F.0D�	�I���_
�u�����|�G�p�P�Cv7X4ki�H8Џ�Ӿ���yi�1tSjv�!�`�(i3��a�Om��)@J����蟯>�������� л��5ߧE4��!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t��&.��8�?9��I�f���ܐ�}�闶P���`�3ޕ s�O;,�	�;g�x���o�˩&���^�``��yJŹI̄�ѭ����V��$�� ��D��)G����x�p�8	�W���
uH��Sy8����a��)9��.o��ְn����4����h�r��~F�iO	���gL��=�H65�������D��%C1��,2�A���ۖ��S�<Ԣ�:��ڂ�KQ�������\F�7��0BA��_�+m�(��k81aJ= 2�6�o8:4�I���c�90@�ٍD+��z�H4l�N��b���Qw�c4~Nr_�mS8<�nE��6�3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�V�һ�d��[0����F��5��܊K�+���w�PjI^�UI0���ԏ�.fOe	aNq�*��!���Q
ŚA���ۖ"'��&އ���lc�ڕ3��t�>�!�(Y�*qA����6\�4�@�� �-j�n
V~$�=���\%��8��GM�v�]��1���U�._�h�5,Wlr�r%)cA/�r�]/2n�����$��@%��>M���b��v݋N������$2ܓ�A֍�a-6�DaR\�^.����c�v�J��sr�l�k]m��^~W���e�G&�A���c�v�J��sr�l�k]m��^~W�����5Lwn�3
�v�v-}�	mpBR9ƭ�����fx'v�ao.\C�k�Y�\�p8�<l�o�>>����I���I�����OeU���(���,�	%���_T���a�aq����i��on
V~$!+���}���gn�=4�4�	���WdM4@�肥�J�O@�s��M���c�v�J��sr�l�k]m��^~W�����5Lwn�3
�v�v-}�	mp��"����I0���ԏ�.fOe	�HlU�!=�����gPh�Qf��o�U/]�i��N�Na����g�6���Q,|��,�ϣ퉧:��oQ�|i��N�Na����g�6���Q,|h���fn�g��]�J*�Rs�08�b(��z�X
3kZ�c¦�.��q��`�L�����gPi�a�sirUë��FWҵ�3�L����e�eV�M�z$��P�!�A˪[	��*3)�����3�L����e�eV�M�z$��P�!�A˪[	�$^J�����fx'v�ao.\C�k�Y�\�p8�<l�o�>>����I���I�����OeU���(�1O,J��I0���ԏ�.fOe	� 	���R�h�Qf��o�U/]�i��N�Na����g�6���Q,|��,�ϣ��19TH��u��)o���r_��m����&�Ko���&�@�}7�q��J��v1a{J�h�µj�!�.M�LYq^���&�@�}7�q��J��v1a{J�h�µj�!�X�:�{���zR���b�5ߧE4��zR���b�5ߧE4��zR���bn��9z�v��k]m��z	�LYE�Ut�\�(2ڭt>��b�'Be���0��_��fx'v�ao.\C�k+M����ǿzR���b��˓#���3�5�I�]�C�x!�H�k��^)������K�+���w��ba!؇/�n�����F��O�n��ݕ^)��٥���F��O����Z���׏�����Mc¦�.���IX0F�M�}�I�Ҡ8jH�G�NJ�;�=����qj5�w�R���y��M�~���,ۚ��7\��.�b�U�[2�a%�Gb�+=tg()��ikp���H����~���B�#g�k��m���f�|�]A1�;���o�vŵ����t�T��?E-h��`f���s�������������]�0�zG��"Όd)��u��a��i��N�Na����g�6���Q,|��,�ϣ��19TH���*?�a�ǫcЉ�M� �,ﯾaϡE䦛1��l��=5;vĹbҼ�P��z(2����^a�nu4Bޗ��jw�	����/�ciJ��Yu��&���E��}�XƤ5_���M���R��ӟ-���J��RQ�1z���IdN�^�%��>M���b��v݋N������$2ܓ�A֍�a-6�Dax�Hr�6w��]W�I))����A�m�(��ʢ
wJ�	�LÆ�b���[Q�܍w�S}�zR���bJ�%Ph�r^m"�OB7A�SW�N����4�P��/ ںW|��6����&�@�}7�q��J��v1a{J�}D7B��#��.M�LYq^���&�@�}7�q��J��v1a{J�}D7B��#�ڮ��(�a)x�?{���x.�Knq��!cI͸I))����A�m�(��C��AF�Р=��'e����&�@�}7�q��J��v1a{J�h�µj�!x������_�n�To�[�C��-���m ޶&�hbvk~�#x/����<	��c��*��G�\�4���gn�=4�4�	���WdM4@�肥�J�O@�s��M���c�v�J��sr�l�k]m��^~W����S��]T�3
�v�v-}�	mp�Fy����I0���ԏ�.fOe	�HlU�!=T۳�͕��~K
eڟ7���&�@�}7�q��J��v1a{J�h�µj�!�.M�LYq^���&�@�}7�q��J��v1a{J�h�µj�!vgrEs�1�g()��ikp���H���y���@�Krw�&�z<a��r�����˓#���W|��6����&�@�}7�q��J��v1a{J�h�µj�!�.M�LYq^���&�@�}7�q��J��v1a{J�h�µj�!���H��ҷ&|���BY��l��=5;N�����O�9�d�L��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$
��.�_�n�To�[�}�~��l�܍w�S}N��-���'���c�v�J��sr�l�k]m��^~W����>q�[��q�)]Q�x��r_��mzf	�$NT�I���I�����OeU���(;)(F�T��̙�R��I���I�����OeU���(h�a��Mg.6�kJ�1��씑�:��KY׏�����Mrw�&�z<a�%3�0:=�O�-v�*�Va�ir�4br��`�s�T�Ο?�R��n}�����H�X��WG ���,�%�Yd�Z��2�m�k]m��z	�LYE�Ut�\����7�P�K�+���w�PjI^�UI0���ԏ�.fOe	��<�����B�R���>_�1�<T�b�'Be���0��_N��	�Ȓ�cЉ�M:��V�_��c�}���Fo|k�LbV���G��׏�����MJ�1���۪	�}a�IX0F�M�W/��WuB=�r��C���,��K���Y�q??�d���&�uU��U���Ep�7�$�rrwȀ���3�L���'s{	�h�v1a{J�h�µj�!W�/�#+*f��3�L����e�eV�M�z$��PЏ)�6!@O�O�'�j3Q�I���I���C1zh�6���Q,|]���#�KF��D1c��I���I�����OeU���(�1Xz����4br�����w���9٠��WJG�r�c �4br��o�*�g���OB@1I�kI���Y/������T��"l�A���ݤV���^'���I���φ��<�6�@a� ��fFMqlg��èVxjzӝ���I(͂X��WG �����ͻ�da=�&./���(�6��N��D�D$���1�?��,�����*ւ$զ-�F��,	���~#G��b�'Be��/�y@�,�Y\�C�x!�H�k��^)]� ���_�hbvk~�#x���D�#3��,�-��L��)܅������!<�C�x!�H�k��^)�c/V��"Y�l��=5;vĹbҼ���#�;�3
�v�v-}�	mpWZD�H� �|,��@��(��X��4��VJΣ8��3�L����e�eV�M�z$��P�!�A˪[	�܆�VwB�3
�v�v-}�	mp�|"�.���3R�e��Ӵ�"�6j��;٬sf.�r� F�3N�V�һ�d��X/�S)�5�;���N���A*g()��ikp���H�����U���+��.ᬵy��+��'�׭)x�?{���x.�Knqvcyt���󑟇���-hbvk~�#x���)kb4��VJΣ8��3�L���'s{	�h�v1a{J�h�µj�!�M��hbD��ڙ�n�ZLN�	���}���x�A���ۖ��1�:��o[�a����c�v�_����J�����&����˶�Ka��m�%�\����*\�9X����[JM�D2\1z���@qP<p�CB|�����J6����"'��l������O05 S�s�l�3
�v�v-}�	mp��"����I0���ԏ�.fOe	j�3A������0i�����I��ďr����.�aq��9��,=O�󑟇���-hbvk~�#x���)kb��Yk���0��H��k$�,�
2�[�i�aSA*���:���:��ά�sEv���2�ę�u'b�'=�(f����Hׇ3
�v�v-}�	mp��"����I0���ԏ�.fOe	j�3A������0i��Y��f������&J�b, ӫ/��m�B�K��1Ҹ�]��0�ȍ�x�>c��w��'o�<���q��q+����>(\�H��/Sg�w��'o����=�ɲ�cz���Ӵ�"�6j��;٬sf.��vd��#۸g()��ikp���H���h�Mۖ��V��h�ӵeo��C��=�d�*�,_�n�To�[�C��-���I����Ɖ�Uʚ7�ܩ�.fOe	p�Qz�XO�9��IM� I0���ԏ�.fOe	`�R��7
ɴ��z�4�	���WdM4@�m�"-G@���T�8ƾ?2�?⨣�~��)�A8�%<}���"'��l����C1zhi�Y
�,��'�PD�����g�Z��3��a���!@�f")u��r��܌;���d��-��!�L�F.	-�L��&PY~�y����o)�T*�c��܍w�S};|>r:w����M��2Ď3��D!��;e��J_�d�@���GS滑����ZLN�	��MdGN����u��XC���}D՛��W;���\�H��/Sg�w��'o�MdGN����W)�x�F[�-6�$�D	T;�i�� ӫ/��mR�MP��G��]�,���;���N�GT&D����a-6�Da
] +S�u�v"h�`�t�2�H?�0��b��Z[�MD�ԱC������gn�=4�4�	���WdM4@�肥�J��eqm����gn�=4�4�	���WdM4@�肥�J�����Z����"~6���aq��H�&l�u�&|���BY��l��=5;N�����O�9�d�L��3R�e��Ӵ�"�6j��;٬sf.�r� F�3NNq�dd:�g()��ikp���H����濫�L�ፎa-6�Dazf	�$NT�I���I�����OeU���(;�~1��_��	�_��:��u���'b�'=�(J�}�֖���p�5�Ѱs��訌��v�8:��˗�a«��fx'v�ao.\C�k�Y�\����pP�h�Qf��3R�e��Ӵ�"�6j��;٬sf.�r� F�3NA�׭�%*b�3R�e��Ӵ�"�6j��;٬sf.�r� F�3N�/%\��jX�m ޶&�hbvk~�#x�%��4�w3t���=�4�04�jfB�R���>_
H�n b�5���c�v�J��sr�l�k]m��n���=�y�e�G&�A���c�v�J��sr�l�k]m��n���=�y�kU�����>��� ӫ/��mt������9�d�L��3R�e��Ӵ�"�6j��;٬sf.�r� F�3N
��.�_�n�To�[�}�~��l�܍w�S}~K
eڟ7���&�@�}7�q��J��v1a{J�}D7B��#� ��JJ��T���pP�$D\��z���gn�=4�4�	���WdM4@��&����˶�eqm����gn�=4�4�	���WdM4@��&����˶:�D5��h7�P�HS|�4�04�jfJ�1����ݾ-/�o|k�Lb#.w^�oG��8��GM�v�]��1âq�t�dh�^V��h�5,Wlr�r%)cA/�r�]/2n��ɲ�cz���Ӵ�"�6j��;٬sf.���Y�m��
ɴ��z�4�	���WdM4@ȁ%B�\�Db��E(�\�H��/Sg�w��'o�9���&aD�4���t]���8����0�J����!�(=�oaJ����2�/��Q��i�<�t~f��X������UGɤ��g�X��9&���K:+>����YxP���2�ę�u'b�'=�([>	�ە����a-6�Da��zb����2�ę�u'b�'=�(xa�s^����o���*ٝ�/�K^b�;��	+�}�&�}�T۳�͕������4~V#�(�>^�l��e�eV�>�3�eZ~�/t����"'��l������O&�4�_�c�}���Fo|k�Lb��@^�11|u='�c�a����gi�Y
�,�LٗH�1�"'��l������O�N�ʶ�L��zĐ��OJ*�Rs�08�b(��J|WQ	��2�b��v݋N�����|�+��)�Kh�4dZ�Ր������aA�(�W[��nn���t�3?r*B�#<�T�R��OO���EH�a���#_/<�I�i��a�z6�&aD�4���t]������o�*����H5��M�S��X���/̥@X�4��@^�11|u='�c�a����gi�Y
�,�LٗH�1�"'��l����C1zhT
�����=�����|$�b#���:>���b�<~ ӫ/��mt������9�d�L�ɲ�cz���ł)w���m�±��m|����>��s��|��袔MUt��!�R�x�ky~K
eڟ7C��(3��7�q��J������-VL�4%�YE:�|u='�c�-��;���_�vԡ3є�,hy�̥͌!���5V����o���*ٝ�/�K^b�;��	+���:��KY�[b%Ɨ�8�%<}���"'��l������O05 S�s�lɲ�cz���ł)w���m�±��m|�b��Č�?��|��袔MUt��!�HlU�!=�5ߧE4��p�-a�D͢bP�63Z�t��Ě����z%�ژ�(�*4��%�#o�]�ʄ�q�����~=&lL�i��D!�0�?�R��n}�����H�X��WG ���f��^��z-�39��X��WG ��W|��6�C��(3���-��w��k]m���.M�LYq^C��(3���-��w��k]m�����H��ҷ�Gr�}��_�n�To�[���9�P�4�K:+>����YxP�B�>��֑xGV�-��\�K�+p���#4�Te͉�XkN��"�&CX��WG ������4~V#�(�>^�l�'s{	�h�����-VLU4���Z��"L?���N��-���'�[�s���_����J����:�4�k��[�s���_����J����C�DF(a�Sc�}���Fo|k�Lbx(�i��/RŻ�&ǥ��bP�63Z�t�5ߧE4��Fr��j�_�Ƭ7~�rG[Pt���匷Q-�dM�V<�'i�*��)�}>���|�X��V�掘�/������-Ӥ�v�79cKAW�������D�v1a{J���Ѫh��*!�Ȃ; ,@�� �5dB��̊�X~��`��OO�����g����1��e��H�P�n����=$$h�8}ջh@�m���Mٙ٣9!pz`  �d{ߥ�L@s3�-�~�.G�ӛ�e��k�J�}�@��h9<���F!+�+$����~���lsه3
�v�v-}�	mp�����W�D<�Gs�B�K��ȅ�"XC}ץE���������J�)��Z+���g��o����>�/���M��2��%�;�aq��k�7� r��ŀ��`�z���xl%����v&5��7.�ǖ��`Y�}q^J=��ڥ����Ⱦ|����?��%�th�{X[�QB����.��/��u�}�e��k�J�B�Q����9<���F!+�+$����Z�8	J#�=9���G�n��<��%m�Y$� 1H��!i��6U(�<";)(F�T�M�{�|Lɥ���dh��B��p��XD<�Gs�B�K��ȅ�"XC}ץE����uB�F8�����J�g���ʥ?�v��7�����Ȕ���|b�}�vy�
�eʣ͜��l�l�A5�[%�$�r�ի�!�)]���}�Wy5nTf��8�i_;�.#x��EHhYOZ㫶��`.,�`�_��Q��R������6U(�<";�~1��_��M�{�|Lɥ���dh��r�f87�&�<om���m-F���TX[�QB����.��/��u�}�e��k�J�B�Q����9<���Fv &~N�gr��Q0e[P!��|����GuDc%^oe�Y4)_5���ʮ�&*����}g]�X�P�(?`����9�/�!nU��K.��QW�4*(�$���W���[�����zޥx�
��J�f'o�~z5=����t�m�՟��HN�2��$cC�Z�_Ԕɺ6�r�>�e`�=�a^�e8�b,7��6~�p�@OM.Ir�b����g������J*�Rs�08�b(��@��C2K�ǽ$�!b����#�GWW�<om��H/�>��=�M����ge���ޒ�z���t]������^�k/^���H> �s�bͦ-(����U�._�[t�Y81�d�@���G�X���.��ġ��,���'
�?��p��6�>�b�WI�F{O؏����:_TqaV���M�{�|Lɥ���dh����50f
V��.ᬵy���Ÿ�`u�V-�*yT��XƤ5_���"~6���aq����i��o%m�Y$� 1��3�a䗉��`.�eV�U��)���Y;e�iK ����)c{y����i�q,?5q�p�'�ˢݱ)"/ǭ0�zG��"Όd)���jz�\=�/��8y�����Ϝ�F���[�4�f,�{_8�Y��=�}�Vݨ��&��M�|�+4K-����)~u4���܂E�g�������(ӈ��� �3�c`�k+Q�h'�Ȝx�5W ��̫(>��o���,l����M?��y��L��Y�_��&7�䬬��_=���z��2�^���6U(�<"j`�RU=�R�wX���L��Y�_��&7��������z��2�^���6U(�<"�lp'^��gR�wX��rw�&�z<a��N� ��M�W8߸��S�Ȍ�w��ڷoy��� k���-�+n̪p��9����~���=���q5�nn��e����;��|B�R��Ρ�U�MMk�R��6�o8:4�I���c�90��B�O>qiI9�o«IX0F�M���H9U5���U�u!��I(͂X��WG ������CU��O؏����:�xH��{as���}�pIɽ�Jz_ꛨg��U-�e>� {�}���my$�N���Uە��g����Ǵ=��!��������LO1	3i�\��׹��t˔R��}K7͍��wAA�Ɓ=<�W�.�P�Զ��ߘ������g�Z��3��a���!@�f")Ut�\�e<�Ia��la��o���1�ź���$��Ly��l�7�wۤ��D��+_���R̕q���s���4���܂�c�eC(�55�k80���렵�!E�Y�G�˱�ߓC娤l��°������R�wX���	G�˂�c�fi�dL��_���/�n>�.-,��Sq'���Jy{���C�|J3J���\&<���2u?r���Y�G�˱�ߓC娤l��3���W
�rw�&�z<aSm�6��`4�04�jf��ܐ�}�|&�xVgY�b��ٞ@[�_zβrE��g�Hb��-�+n̪��0čK����uwn��e8�b,�9�@�Xc�v����O؏����:ջ�F=�|�!��AHFu�ﶲ��Cҷ��e�2�^���6U(�<"�lp'^��gR�wX��O���M3X*��L1�]RD§B �����+&go#��S���*�7G�zV��� N٣�RD§B ���`y����	0��E�ǖ��`Y�R}��کe��k�J��ֽ�\���� ��pE����CѼ���ߙ4�� �#��S���*A��� 2����k����i�rd��������c�eC(�5_��&7���7M=�L�f~��DV��O8�#7S������6U(�<"�˨a	e�!�6UVoā"�z��h,��J�`cL�6�9x�cx�Pu9� ȫ^��t7!CX~�
)����Ҥk����x��'[W����E !+��=H~3�A�Â�v��c�/�	6������1�R+-h]��.�{+��f���i\�H��/Sg�w��'o�?S�B3�<X��kRCլ�����`�� a⣃_B�~ޙ����fQ����2I��� �'d��0�˽�}ޡ[�aBa �k<�]X��˒�Û���G�'�����{��-Q�=U�KO���d��s���E�n���
Ո�C�hk��Y��A�m�(�RB���
��\�� ӫ/��m2���K��֌I�<�������|I�ݱHه��;��|B�2����&::��n[I?��8y����e��s�ZI��RhF��j���W��׹��t��h�	�Ȟ�����Ao�2�P�4x`�1)W�w��fD	���%�� U2�h=c�ن���8+c�WT�D�3�=�g��������s.'�����'�� �4&OKyl� mr�m�e*4��O*%΢Ӟe�a�f+(��at,�9�i"�e8�b,��fC��rJ[�x�I�"����Je��v��YN
��)e��*-�3Y`���$� ���U� ��V�I�Q`���$���^��y6�T���1��豁��P����S����Gd�^��z\B�IX0F�MV�ҁGG��ABk@�`���φ��<�6���n�4��������]�0�zG��"Όd)��u��a��i��N�Na����g�6���Q,|�b��暴�ܴ8`���r%��ɷy�8��O|E�g�������=����z�����y��gn�=4�4�	���WdM4@��&����˶1X�iRd��D�����X���*"��Zʊӽ����K7͍���\C�
<rg����Ǵ=O�W;D�1X�iRd��D�����X���*"��Zʊӽ����K7͍��wAA�Ɓ=<�W�.�P�Զ��ߘ������g�Z��3��a���!@�f")�4v!4���=�O�-v�*_�mS8<�n�$�|�K��3R�e��Ӵ�"�6j��;٬sf.�
�DB�%�$�nR��ړC娤l����pQ�q��!W�	�_��:��u���'b�'=�(J�}�֖�â"���O�׹��t��`�J9�������S���v�+��gn�=4�4�	���WdM4@��&����˶1X�iRd��D�����X���*"��Zʊӽ�����3R�e��Ӵ�"�6j��;٬sf.�r� F�3N�f�uj��f�C娤l����pQ�|f>����B��eS ��"��������LO1���q5�n-�@�4ڧ%�fL[���o���FO�W;D�t��S�D�����X���*"��Z���Q3��p�-a�D͢fU�9�׏�����MFi��|����A�;��=�#�5n����%�;��|B���~���}0��u�X3�����ۺ����� ���Jx�y�Zgl�.�����>Z[t���{�ag0Rm� �[ >�3 ��V�I��`��ٞ�R̕q���'O�����Z���4�+Mi�C�G����]'\gWg��	�Z�kfc�Q�bc�+:Fa�7���W"�P�K��q��[@����U�u!��I(͂X��WG ����rzj�#��v1a{J�|����$/�pX��� xh�Ɛg)x�D�����X�0������my$�N��w�ci��ˇpPo��zX�C���������C��֑xGV�eU���(n��_l)�t	3i�\��׹��t˔R��}K7͍���\C�
<r����4~V��3�L���'s{	�h�v1a{J���>	�`�`��ٞ�R̕q������鷂�nF���W�_te$�J�� ,��8y����+f�8�ï,��Sq'�@8�Qq���z���nF���<�W�.�P��c3�
_,vF���sݐ��,���$:N��@�1�˓����Uh1�b_X�XV�b�z'hۉ)��R����\�G�����dc�@c�����hX��WG ��������M���LQ�/8qߟ��l���\�.�۟�n�O��Ե�	3i�\��׹��t�M��|S�/���[�4�f,/��U���JVX
���$:N�t%��zxa(􆿳�e�&���6��ڭ��*���!��|�Ɛg)x�D�����X��Q��Y��O\���򙷉8y����*S����,��Sq'�����f�՜�T�\ ��z�X
3kZ��*?�a�ǫcЉ�M��7�ጰ/y�搲)���$:N�8.����6��DKY���k]m��v��z_�Ŭ>�Y�G�˱�ߓC娤l��3���W
�~K
eڟ7���&�@�}�-��w��k]m���%�8��>�y�搲)���$:N�8.����6W�/�#+*f��3�L���'s{	�h�v1a{J��8���-R��`��ٞ�R̕q��]I�3�z�X
3kZ�X�C���������C��֑xGV�eU���(�˃��'�	3i�\��׹��t˔R��}�3R�e��ł)w���m�±��m|J�}�֖���6Ř��%Y�G�˱�ߓC娤l��3���W
�p�-a�D͢q��`�L�5ߧE4���������~�LqJ��.
u�Tг��S�?�d���&�a{�(%��r%t�PDa]6j�"HsF�prB/�*@�/뱍G���6υŽdkYF����o�~��V(����\��K��G��*�/5�si鏈wƠ���z�Ig��mQ3��T�2�1��o2"35�&P����NJ�q)�K����ȑ�z�P���(fw������C4�֮��k����H�V�n8�A�A�/������Z��Ջ\{ف(�7���`�z����k!�\Z��K��qb	��G���Q��x�/�����y���|���������S�_
�u:�_q�pWK�+���w�1��Y���;����;^�6#9>���@]�E�i�m}66j�"Hs1��i�����s����aT��3G?�d���&����AW �[�p�*v��)����o�>|/���H:>�� ���Jx�y�Zgl��>����C;��|B���S#���회�h�#5ġ��x���u�Y�KG�ξ���e�J�Pn\�pD��ZOU;��|B���S#����b�'Be������>���$���gE�s@�j����tL���.���k]m������ˤoP;��|Bɨ ���`��s�`DVB���_V�|W�w��fD6S��^[�p�*v���q�	��c�d�e?��9�V��r��N[ m�N�P�ϫ)+��'{����O�L�0��i=B'�{3�.��"�l�j����+�=�z˥���#���F�&� &��(���H�V�+R��}y^���L�D�d��2=��h��IX0F�MV�ҁGG%4vkz���յ[+8��r$ɓǃl[�Ƶ�1tSjv����8�2��w��kf�Q������(ӈ��Z��&61@���rahv���7�R � ��|��5��9	v�(�$�T�z>�Z�n`J��@CJ?\,Qö5��4QI�T`����`��HM#�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�����㱼R�o��ob$fAԢ�a\蟟Q��ǺΕR��ӟ-�q�x�~<��w���	�e���(��6@g7����U�._�3
�v�v-}�	mp�JN�7��u��r��;�jmT�#�T�n��a�j��	~�<om����J��RQH�RtV�^��{$@d�̟�1��{!0g|���#�=3!�`�(i31���~!�`�(i3�T�n��aγ �,ﯾa�ݚ�Н�$f��_Ub���r��������_�N5�Hɫ˨Â��P�<om����J��RQH�RtV�^��{$@d�"����DZ�NU�d�@���GCq;�~����}Dq�f��	��x��ݚ�Н��'.�T��ol��Ә�|ƀ��K_����d�bfĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹���	Z�;�|��L�D�d� {�'#������,�ǰ	M,��rER��S�p�����(�t���pA2wKaC��=}'t<��ġ��,Q17�b����#g�k��ö5��4Q�]�p� �)R�G�׵12�mj� ��JJ��T����,�ǰTm�v��G��d�@���G%fE�g�=�&��q>�<�'���I����� ���JH����8����F)�~����H�V�n8�A�A�y���6���#¯��TG6�o8:4�I���c�90B3v�A����èV\���F�`yx�>�+X�M?��y�!�`�(i3�4br��n��>�my$�N���Uە��g����Ǵ=�a�D��<F��� ��f�{_8�Y��=�}�VݨuN�wAB��O���&z� :�:���^�{�&�R��\RU\Dn��c�L�{�t�� �?�;$^7E�g�������(ӈ��-�G�~�h-:���h��T�٥��T}�a�mC�0��\RU\DnscX{�X!,	�)��&ghRV��R���P�|T����{7�H����8���O�υ���YN
��)e#j�o����:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3�I��� g�����Օ��qvdЧ^{�jMdGN���!�`�(i3%Q�[�J����˦G��4br��6 y2��R�՝� s�#���k$ �B�'��a����aGl���nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN!�`�(i3]���-_!Q���ŴIh�5,Wlr�r%)cA/�r�]/2�ݚ�Н��ߎ ��E�VTҝD!u���o���F������}Dq�f��	��x��ݚ�Н��ߎ ��E�VTҝD!u��nF���<�W�.�P�	��
�Q�}���%>�rG4�04�jf(��Vb�h�^V��_�mS8<�nvE7�MW���㱼R�~=&lL�iX���\@j?�R��n}�����H�X��WG ���	G�˂�c�fi�d5X�nd����YN
��)e�
��9�ܺsl/=��"L?���M��ZLh-S���%��V�c��݂�nF���<�W�.�P��c3�J�1��씑�:��KY׏�����M�; T����%�_�n��1q�JOG��Hb��a-6�DaM-��&���������Ц���Օ��qvdЧ^{�jMdGN���M��ZLh-S���%����g���hZ���o���Fq@L����?Y��Yf�>je`��@d:�����{~�
\za$Ad�*8Җ�N�>f5�� b�z'hۉ)��R���p�-a�D͢q��`�Lx(�i��/R�ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��׏����y���6����8��`������,�ǰ	M,��rERu!/��"��H�6 ��Y%ɫTKA2wKaC�(fw���'�̗������k2m�;��|BkCD��9'�̟�1OW�fL�
\za$Ad�e�h�`^Drp�叧w�kkr�i�<�j�&�E�g�������(ӈ����L��c,S���%����g���hZx����E2b�z'hۉ)��d�7�qĜ���,�ǰTm�v��G��4br��]E�'�f��ja5=��)Q��U��)���Y;e�iK!���d.���8-|�D���"sS<�0�zG�������&G0׊�E�)�̟�1�h�N#�Ǐ.qѐ��_O�4��"�V�w_��Ǹ���)/�~�T���]'�^��������F�e%��5�J\��+ʛ����{_8�Y��=�}�Vݨ!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^e<�Ia��la��o���H�RtV�^��i�:�3>�XƤ5_���M���R��ӟ-��濫�L�ᙣWv
*T�>k�N��^��hJL��;���N0�!5R�Ut�\��H��Pk	l�
@\ه3
�v�v-}�	mp5���%�+� h�ҩ��wӨj]h��Z�8	J#�>�8� \p�r~�h��ݚ�Н���w�w:�݆TO��My����iI�^օ?D^��!�`�(i3�5ߧE4��!�`�(i3�5ߧE4���D�$0��4br���qP�V>t'�̗������^ā�Ӱ1tSjv�����l�����r4����$A�S��b��v݋N������$2ܓ�A�� h�ҩ��>=���#�-6�$�D7���s�a'���c�e�C-��[
�:qEp�[b%Ɨ���:��Y1�s �n#;8���'�PD����%>�rGO�D mWN���%>�rG4�04�jfx(�i��/R#.w^�oG��8��GMӫz�Ζ�"���7������Lh�5,Wlr�r%)cAH�Ћ�r�\Bk�	��^� �S������2=�>c,����{���3��;A,D�
���kC/��E������GI��	r0�'�Y~�y�����?�J��܍w�S}�W)�x�F[�-6�$�DK�(+�`W��,8����;A3�@���Y֍�a-6�Da>f��8�D�u��u���)������ɛ�?өT۳�͕��u�޽�vUMa0��#��������"��=�<�^p�-a�D͢q��`�L��˓#���9�x?4:��-6�$�D;�,th�5�۪o�y)	�'��ɡ����4$E�-M�O��~��W)�x�F[�-6�$�D;�,th�5�۪o�y)	�'��ɡ��y�A�?�-M�O��~���.�2��0tNF5��q���v�{%��v��>je`��@d:�����{~6�!˓C���I�Au����V�hdW��Hp9���5ߧE4��p�-a�D͢bP�63Z�t��Ě����z%�ژ�(�*4��%�G��Hb�3�� �f���r4���(���q����M��2�B���l�2��Fm�ӫz�Ζ�XƤ5_���M���R��ӟ-��濫�L�ፎa-6�Da�N�]�B���vE�fc��57�Mv!���xFhMV(@|΁-6�$�D?b{yt��>�۪o�y)	�'��ɡ��x�s�?U�H�-��pQ��e��>��Օ��qvdЧ^{�j��:����
�hf���CK)�yynmg�ibZ+���g���+���8�׏�����M�4O/3�L�3B�\GJ�8;��w�h��Jc'�yK�w��g��U-�e�՘�L3�CK)�yynmg�ib��6@�������΁In*42�����`y����;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6���ޡ�m���Y�$����!Oe�Ǹ���)/�~�T���]�^0���7CK)�yynmg�ib��6@�������΁In�D�;F�)2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�S*�"�=3�Ҥ�P�X��������3R��kѶ���� ��&��h�?i�H��}��?<����G&�;���� ����}p閭3u��N�,?��΃���]�X�ֻla�oZx�i�xx�j�甯�[���pФq�Ǒ)''��m�9X��W��� �_%B71Ձ"�Ĭt�'�ǅ@s�-6��P�%Ae!�`�(i3<�6�Q=������Kd���{J��&�~�����t�tS�SaqZXr&ߜ�ۛ�&��#����^wO�L�=F.�,��J�X�:zJy=~�*���-�������ó�$R��2����C��P��I2��0�е�5<���3B�Hj7h~S܄=�չ���1�]�V�#0ݱ���`�~�26��\�)�!�L��I 1��6�pa�Y%�^��g�ZS^���\�}����P���LȬ@VYBWh)b�����k-�c�����M�~���i��lH�I���[�?O;��c���X�ʛ_��@ a⣃_B�=�WK=ZȞ���]dF!�O+�|fc��57�չ���1p�z��.gC��	����Ow���]'\gWg��	�Z�kfc?�#	*]]�(&�L�xjzӝ���I(͂��-����r�VU���N�\�]
��s�G��38����]dF!�O+�|x������a4���܂E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*_�mS8<�n�ݚ�Н�JnFݲ��s�5�>U�m�j*��{�%L_��f�����,���R�e�0����[�4�f,�'�f��P���U+��_���|��5�>U�m����9gUS�|#9���
�:qEp�;�P�t�5fĉ>99��A0ok�׹�R��l��+ݭ�~r}�!��sc���!���{�'�f��P���U+��_���|��5�>U�m�����ڗ��V�=K'sR;��|BѪÝ���/����u��u:u����<�Zz�a�h�5,Wlr�r%)cAQ17�b�����d���!it�td���5�kv޶Gl8��?|�,�e��0�U+�qbp@�s5]N�uA�ۥ�Y�m�չ���1�]����7����0�;�Fi��q�>Ш��+��t,�� .6�o8:4�I���c�90B3v�A��ʃK�,��`U��B��-����A�;�����\�5ｵ����<�6�Q=�r$ɓǃl[�Ƶ�1tSjv��� л�Sm�f�e��N�eM�#��}Dq�f���b��~�F�KD�Vr[/}>5��0�B� �b�в��y��lD��KJP#�'����u��r��<�6�Q=�dOP�m�(�Ha׮�#K���~N|O`�� \)0��l!���O�D mWN��\ Nh�;�P�t�50��l!���߸��S�Ȍ����[7Y'��k��F$�kj���;�Q�s��'G�+p�Dʾ��6�o8:4�I���c�90B3v�A��ʃK�,��`U��B��-ն'�U;|�u}D��� q��j�J^���{���#�0�zG�������&G���y��lD(�D �6��Z�H��q�e��0�U+�qbp@�<�6�Q=*qA����6\�4�@�� �-j�1tSjv��� л�e<�Ia��lb~*��s�닓.�`�3+,w	�Af̓@?5�a��ToEn�A���ۖ"'��&އ8�fk!�`�(i3T��a⨯�d��+��2VP��Ѣ�ʒN�ċ���y��lD&[�x�R�"��}Dq�f���&.��8�}Q�sd��]� )�+����򙷜�9���w'-���JN-Y&yo�q����,�ǰ����adp��e���W�~��$g龙]C�1�ɕ7'K[�� ���JH����8����F)�~����H�V�r�Z����Sm�f�e8�1ޞ��&e[u�;0�2����k�����#�K�v,���cL�Ec'�\Y-φ��<�6�@a� ��fFMqlg�2N��n�O#H��EkנaA<���XP��Ȩ���[1�`���φ��<�6��o�.�u:u����<Srƫp��xjzӝ���I(͂��-����<�6�Q=����P%��v��!�`�(i35���u�L�����y�]�"��^9r�`�	��'DV���b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^hs�����F;p�	1x�a��2'���Xw�j�7�����P�|T���;���%�����T�`��9d��Ί_����ݚ�Н�|�au�(Z���Ma�B�#y�D�5�S�`�	�ӛ�i��.�mJ�0�6�!�`�(i36��J��c��Yu��rP&��dGL� ���8#�Y~�y����o)�T*�c���-/a8!�`�(i3pi�NWHC�ۥ�Y�m���NM���!�`�(i3-6���[��<�p��Ar�8w�B
�:qEp�gdq�_x����Yzw��(4G��>��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3�$VǽO���!���{��b+}y[!�`�(i3��NƥNoz��KUq!�`�(i3�����!�`�(i3pi�NWHC�ۥ�Y�m�չ���1�]����7���V�� -+;X���W���b�0����%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ī:f����p=�3Yj>��q`@D�[�Wx����'G�+p�Dʾ��6�o8:4�I���c�90B3v�A��ʃK�,��`U��B��-ն'�U;|�u}D��� q��j�J^���{���#�0�zG�������&G���y��lD(�D �6��Z�H��q�e��0�U+�qbp@�<�6�Q=*qA����6\�4�@�� �-j�1tSjv��� л�e<�Ia��lb~*��s�닓.�`�3p��2�H����y��lD�l"�C��XƤ5_��,\���*s-�e�2>J*�Rs�08�b(����T�\yb�����Z>��A�$�|���y��lD�p5j\"���XƤ5_��,\���q���7?�R��n��/�����{N`�/~��խdp��;�{��!�`�(i3���E?����׽���H+�����Dv�/"sB!�`�(i3��&.��8�F�S�1 �烉s)�v�bP�63Z�t�u��I��g��ޏ��ʦ�X⦫w'-���J��;_��8W�w��fD�]C�1��l�Gm%61c¦�.���&T�ͪ͌�#}�{�Ɠ%�ބ@j.�0S��U��)���Y;e�iK!���d.���+�^n=\f�5>��؊ګ�$������r$ɓǃl[�Ƶ�1tSjv��r���h�0�I����~u/��kOT���q�D��1���~��/��kOT*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��N��W��pp�N1U�Xr&ߜ��[~5�{ �q��]����!'PiY�����$��%����ht��p���_���{$f��_Ub�d,��B���ʬw�S���[�Z8&�Ut�\�.�V4q����`�_ 4��;�P�t�5$f��_Ub���uQL+��φ��<�6��9;��ˉ�z~Z�����DZ���I����~up�@OM.Ir����|��6VAtD�/��,�z��g�չ�Ad��x�`�8�G�MTb7-�xc�!{p85v{��lw	S���p%��rװ�p>�"Y\m���DZ��%j_H�ˉ}�@��h� �4&OKy��mh���|�+4K-��T���x2���Ic��AȂ�o�+��5c�u��EeL�V�l��(������}�@��'	�?��[��羹��˙Ǧ�kN5�[՚1Dq��P�<
�[�H���,�'�QDn4��F�(=0��L�r:b�Xϋ?@����sr��A$�P������5d�����Ě���`���φ��<�6�2VP��Ѣ�eʵv|�AәG?��S�0�zG�������&G,���)����}�a�E�Rq���my$�N��o�/���;:Ha��VKk+Q�h'�Ȝx�5W ��̫(�y����A�����Yu�������&G,���)[�л���7Cw�Hm��ոA2t\��,���)���F��O�C#/<���q���F��O���>1Y�$�)�vxV�/e�,�6������P$��Rli����DZ������и;2z��
�@h�5,Wlr�r%)cA��z>9�R��d���!i��D��J�Z�Rj�7�O�e�^E�xa�/ݺ;��|B=y���SS���Q�>�c��)&cm:a(#�ߋ�-�ct�����N*��ј�Օ��qvdЧ^{�jmWᅫw�5�O�%E#P�j؋�������\��]8��	���#�z��%]'\gWg��	�Z�kfc69�#��r���+�^n=\f�5>����Db^<�..�4��<qs��ȓM�Me��=�1��*�
�I(͂��-����<�6�Q=͜��!?@K�q9+t�}�ݚ�Н���Wh�7��2�b=��'DV���b�z'hۉ)��d�7�qĝ�\ Nhk+Q�h'�Ȝx�5W ��̫(� h�ҩγpo守�u�,l����M?��y�!�`�(i3�q�	��c�nz������4�	��E${5j=��!�`�(i3yh� k��4c�!{p85v{��lw	bo N��7�0��l!���O�D mWN��\ Nh�;�P�t�50��l!���߸��S�Ȍ��7���9��e���W�-��ǿ�/��>1Y�V��	��y���x.0 �ιf���M>�����'�=�O�#��iG�taͲaԿ	�Kހ���|�����w?����N����M�\�������
߹��B�φ��<�6�@a� ��fFMqlg8����z�:Fa�7������A����ᳮ�TȓM�Me��=�1��*�
�I(͂��-����<�6�Q=��Q7lY��)P<�ܓ�Y�� л�����g�Z��3��a���!@�f")u��r��;�E����=�O�-v�*_�mS8<�n"�"+U��ݚ�Н�@20߀���c��qVw���%���RAԢ�a\�h��w�{�_��sV�����נ2<�i����)�Sq�l q��j�J^߇�\���*C������ݦ�4����_
�u� خ�^�L˜�,�p���(��6fM�N$r4���1��'��1tSjv����y��lD�;4<�Xݓ�
���T�A�m��y���|e"0��l!���O�D mWN��\ Nh�;�P�t�50��l!���߸��S�Ȍ�"�pӺ^$R��X鷴QW�w��fDT��T�^���h�.xY���ҪQ١Ӿ�$Ջ������U��)���Y;e�iK!���d.0}}��*ꅺS�J\7���z�G�	S�uimK������t5��IM�Ex�>�+X�M?��y�<�6�Q=Q١Ӿ�$/s�1��pE�g�������(ӈ���m�r����@20߀�Y�)�}��EXs70��nF���<�W�.�P�	��
�Q�}��b��~�F�KD�Vr[/}>5��0�B� �b�Ю� л�e<�Ia��la��o���H�RtV�^R���Xc���*�Աߛ+����O��n!%����no;�M#�vzR5�<a��o���H�RtV�^�k���n�9I��@������˦G�R�c4!`ob.�Y�2W>������0��l!���O�D mWN<�6�Q=>��:J�E�<����i"���W�G��!�9Ƞ�������-ќvP�����e��Օ��qvdЧ^{�j�Q;���2� ӫ/��m��?�4D+M���!��� h�ҩή� л�������k��O?���Q�lՖ̮��zՠ�*�S5 ��ݚ�Н���A✵0�ݚ�Н�@20߀�Y�)�}��EXs70��nF���<�W�.�P�	��
�Q�}��\ Nh�;�P�t�5�� л��5ߧE4�흔\ Nh�;�P�t�5烉s)�v��IX0F�MR�c4!`��]��R��M�3e0�g�<����i"��@#('�cH1��<9Oy��]#�0D�	�I���_
�u�_C�7�2������}0n�V2���]#��t�ѕ1��ŦLJ
1H�
!�`�(i3!�`�(i3پ[���-.�y�� #� �,W��-��h��ڥ����ȾY�)�}��EXs7097��EN�y�JB���PY~�y������̡99��: ��ao.\C�k�$���4z��K��zd���|�b��խd�g��;��_���`!�`�(i3}Y;�jn��n��fT�x�:��#�9�Q�f���U�<rM�W�G��!?�d���&���X�իZV�ط�aFmғO�4} ��$�,���n`5�fK�\w��0]����v�E���a�e56<�:�-22�v���+�J���q���U�C#/<���qHe�-�c^Xp�ђ��E����FZ鎬����A��:6])��[��x+%��B@��������/s9�d�٣��>����C�V�ط�aFmғO�4}`L����D:�n`5�fK�\w��0]����v�E���a�e56<��f��E���$ r@{�q���U�C#/<���qHe�-�c��d��]�Q�}J�AZ鎬�������(����F�dHw(��ES���v�8:ۛ@W:���#���FӪ�c�g<�g��U-�e�,���6+�
_g��c�׺8|MW���0o�_o�x�]�V����6��g�Q�q>x׵ �H���i��>�`ʃK�,��`C#/<���q���K1�dѤЭ���ȓM�Me�����{$Z:hx��G��!�`�(i3�NYV�z\+��R�4.����P}�=l�q�������g2���j��M�Mb�:u�w�vG�q�:�&����#|�1�0j�� л��#�l+��B@
��B��+ H	�=��G���v�8:ۛ@W:���#���Ff���'��ݚ�Н��u�qGDnK�]_!C6%K�pıy3�֩�U2P
�{���ݚ�Н��D���R]��ֈS�&I!�`�(i3�Y�M����j��ts���k�+9=�k���n��L�f�\c`���6	D��&8�,�/7����hbvk~�#x ��M��.ᬵy�෺�8�ml<�6�Q=.ӗ�r�(Z+�,�~�7!�`�(i3k S���zǣ©���s�f�I�S�9;/���!�`�(i3-���j_�ܘP{ǣ©���s�f�I�i�	��_�V!�`�(i3-��w¹��<d�,��L�����y��lDu�6/m�Xc]��E���!�`�(i3Q)��Zl�z��SR:g()��ikp���H������7Pr��ġ��,�a��OY��l�+�7#�	�_:iO�A��*/�|��&8�,�"��Z�Z!�`�(i335ݚ�ܨzރ;�{��C�{��M���ဍ��g2���2�9�ԁ���T!�`�(i3�&8�,�3F�蕌ge���y��lD��/?'�M�4�:a��4@Q�/�!�`�(i3:@J/�R�!�`�(i3�$�~c/kx��D(޲��y��lD�b2D��y%�&8�,������	�;�ݚ�Н���^W��k�Q�#<4^�>N0Θ��ݚ�Н��׉8x�)�{� �"czZ������=��e��!�`�(i3Cݮ2���!�`�(i37�_M��f�?ǉ�=񔿄�aB6Э~���VS��I����nX�8j
Jt��)���2�9�xD�̯ƭU��/ӳx��d��]�Q�<�ry^��gΜ��[�����/s98�$��`��7dh�?f�?ǉ�=񔿄�aB6R���e�D�
�~��\��f��E��Ⱦʤ ���� л�)�{� �"�X;p`���2�b=��<�ry^���l��oC�ʪ%��18�$��`��UB�L5wG�!�`�(i3�5��t�e:F�|���m�R�<<�U ,��rQ�VX%����-䤔���8C#/<���q�B�+2�^����W�
L$�c!�`�(i3�e]�#�?�-��w���i��.@B��8C�{�N똴ak�J�a$�Y �t/�(�P���͵��B@���؊N#(K�DJ��-�|,���Ti�w��V����f�z��SR:g()��ikp���H������7Pr��ġ��,�ԙ\���+�@ϕ�@20߀��9]��j�W>l��? Ah�*h,ChW+x⣗�C��ҷ�㗼�?�S���J8����E^��o۪��5/:�� �|������ᳮ�T���t�T��?E-h��`f���s�c�n��X�`���φ��<�6���iE,�p@٢�ԡ�p5��IM�Ex�>�+X�M?��y�!�`�(i3�>8u]�ZL�q9+t�}ȓM�Me���`6X���dc�@c�����h��-����<�6�Q=:
��x�{�\��N�Ś�-����!�`�(i3�>8u]�ZL�	��*��7�*�OH��T7��v��w�K�b��2W hbvk~�#x ��M��.ᬵy��k�t��8*��}Dq�f���Qѳ$G��A0ok��0��l!���O�D mWN��Qѳ$G�φ��<�6���iE,�pzf����ҟU�	Y�����Vvq���i�F�5�j�))�9�X��52�V�e�1�^��hJL��;���N���,'ѧ��"�oi��|��'~'{w#/ B!�`�(i3�eeN� �c�ˆ�A��6j�"Hsi�ŷ ��R�t��-��'��*�-�b�+�