��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�"� r��������:N<��;���Z��4d��{�
��|��Ȋ)zo1���á-�w~��d�������mo�����(����5�a���V��$.:&R�nU���T���딣0&_���X0���2|	p��rw@	@us��n��/�FI���O8�yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|�(����5�a���V��$.:&R�nU���T�����\�4�slom��Q�N�5�%W0�ր� !�zA>(!�o@���q�&2�Z���8fw��[#M����4L"���ې����~I���&���M�|(Q\��(��~��I(K�b	+��~ķDh�D.�1o�����.��:o(~'�@
��,:�Y�ͩ�,�~�B[��Th_&^�� �T�9�Y��6��X ����W)d�H��K��Ap���`"�E+�-_���^*s&QL���BPJ�%�9
Xߞ���������b֡�0��RL�a)'r�Ӟh� ���G�/9{�d���D
���PJ�\�����A�p
˽0?�.���*��� 9ٞM���]��8����t2�}G	p��#}�{�Sc-@G	>��RL�a)��F>x���,�%���pY�� e��x-����l�;H������K#Q�����1�%1�����:�
�~�K�K^Gc7/��#j��;�i1�璠�J�*��f�I��r�O��C��0���۞�^��u�?�L���zZ�Y���;H������K#Q�����1�%1���
�׺R}	C���`'�t?��<6���'�t��,l����k�8���҆�|n��T�{ ��ʥB�2��;��u���^G`J�Й�m��/K5r��!����%�[[e���|���>�
� �AH�*��.�T�{ ��ʥf�nm��mHG���i�P�Gy#����*��jr�4��X	�ƒ��c�w�A��P
T�]���X����PIIN��d�=o����"���	x]̕%�h�Gqc�J�M=
�ٽi"���g�aa�y���bAg�
d�m��+����o5��6V�|��f$ui�V�3ޕ�L��՛�;��4�W�]�a5��6V�|X40��7��XݓAA����~�9�؇�M.9$o��݉�X��R��
�A�`5��\�4�si�W���Y��݅ 00b�������x�o@���q�&ϖe��!���q�L���Q����m�!=�y����h�}���Hے�8Y�&�\�M�C�вC��J�/�_?�hbHp|����#�n�%@ܣ���m2�5�A�E'���M�Պ�s{�tA�~�u��,6o�-��ΐ�?��A�}n���t�o "�xCo9�Z�.�"�K����	x]�G�Lm=�b�7��Mv�9]Sh��3a��$����aa�y����>�u��8#t����nr�O��C��0����"g�����I��s���1�#���Z��\�����Og����n�&\�ƺ���m�!=�y����h�})6D�T��8Y�&�\���
���;Ppo�6�$�PT8��Ì{����V3��p��b��g�|h�03�
� �AH�*��.㤚{y�ڵ�o!f��L_!�pN��i�P�GyϪ+2�Ľ��3rn{����V���	x]�<���e��8�t�~��,�O�W��s�!5�S��H���)��������ҥ{E�?HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�}�Z���ik2)�
}wʭU&H�1��8�h7H�u�ÍeRuw�C?3d,f$�7Q0�"<�F�ٴB�I�SbW9�v�H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3����M�]��7������@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I���ť1k�`d��q�G�+��T��Rc1"�>_�q��.����_42K�,\ަ�It�k\,آ(��7�j2����OtB!�`�(i3jݭ�F�����&]�+�Q��F���x.�Knq������E����F�Z�>)��<H�-��*����Kp&�@���k��!�`�(i3�����5	��{�OF8<z,Ҽ&��6p%�;>4�Rc��ٕ)����i3<�f�D���X���`)馢䃒����Q��K�����!�`�(i37�ܥ��2����*����i��>�`� �@"#��
}oX�4(���k�;�2M�W�Ặ��Ϊ��p8/��e>����Cx�;�x�[�л���7"�,�>E����-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0</���/�u��(�
t��Y�{'%s��.|Z���I7��-5��6��	���`y����*#�m z����Z��o�����
L'���Xw�j�7����w�K����+��dЧ^{�j����#oM|#9���Q3S�����o5��8�TD���rs�i���`�M�	=̞��>���I�Ūe�ǩ"�4s2��ԜF��g.�~R�a(􆿳�ټ*w2�56
���&~^)�E����F��j��\w��0]��b~y� �"�,�>E����-��%Mό���.�Ɏ�#���?\a��4��(�
t�ژq���U�,XG�wz#�9
4�٩�����
L'���Xw�6�:v/l����Sv�ј�"��Z鎬���������o�	�7��r�=N�By3��<�]�!����M[��Ǣ���ꀍ�����5	���]���>����C���"����Y%T��BPe.��xu	�*�QN����q�1Ig�I�?g�f%��h,�qc��[!V���g�uE�EYZ/�矘��-n��I�?g�f%��h,�qc��[�ԏȣ�p�m~|��#&7���Fn����*�X, ���3�ҺMC�^�.�]!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3"�,�>E����]���J���S�<Ԣ�7Z�:1�\mdЧ^{�j`K�=���b�5����`K`�p��'v��a\Y����[7�d|���f���T,!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�;C@�����R���p,��s�p���\�� ��˽��r7ޚY㮭�����'��(��Ja�xZ��j�
�iB{�Z�_��?� Zh�RG�p�P�"i<,��1��yM�׶��	��:�g��U-�eܣ�'>�!��_
�ubF^�[Jh��S�<Ԣ�7Z�:1�\mdЧ^{�j��t�Ǌ��^̽1��R��ӟ-�D�s�A6�&-���x�d�g��ǚ�9�"�5�ʐ��$���Z��oGM�о٫�(�UtW�*X\[$Q��
�̞��>���ԜF����am�Za(􆿳���2����.���;��\u-/���y�8��C"��y��Fp����f���,(���B���ި����x�3�Aga(􆿳�ټ*w2�56�����bp�g� �-��$�K��{Z��rs�i���`�M�	=̞��>���ԜF�����`���W�L�sQ������f���[��R|#9���b!��u��5?�&P-��eS(�e�f���,(���B��ɓ�~Ҡ	��[�)�D#���ߔk�V\�5��|�~�R�wX��}�
�?����D)����lJ��튝�b�Bϱ���w�K����+��dЧ^{�j$��XCp=8�b(��;3��o�r��`y����@����gGT���/ �o�2����Z鎬�������(����F�dHZ�F�\Ȳ�r�r%)cA�%�\B�����x.�Knq�RC�)pb�8���/����,D�6Æ��U���E��8P"G�wk�١��	;q,6KX�#���x.�Knqd��^��R��ӟ-��͗/m*� ��`y���h}Nw����ϣ%�ᄷh��;�y��Fp����ANʂ�g��U-�e,%�0g��ո��U�M��__���Lec�}���AԢ�a\�/��A����d�a�4$�b!��u፥����A_�͸ޫ�(�n`5�fK�\w��0]b!��u���v� 8�e���b��n`5�fK�\w��0]b!��u�L�Y}śT�!�`�(i3�n`5�fK�\w��0]b!��u፨b�e��`!�`�(i3�n`5�fK�\w��0]b!��u�/N2~-��x�f7﹏�n`5�fK�\w��0]b!��u፣I��m�]�e���b��n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��uፕ_�4����	�Qx�d�n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u�l! ʟ{�b���0���n`5�fK��0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��uፍkv޶Gl���m\g��� L�>�0z�cULd�g>57<�C�u)�6�3A�)OqЈ�&��g3�g��U-�e�j���s�Bd����t���A��'�����ޙ��E����F��1tǚOqB���یHKz�Q��q��3���5�O�%E#P{y����M�V<�'�����~?�ni��Lt���hm�(��k8�P��3���o��_�Rv�䩲$���dS@Ɵ�od�G}%����3f3_�n^�	$m��M[K{�����s#��H����Qw�c4~Nr_�mS8<�n!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+Q3S�����p��8��{_8�Y��=�}�Vݨž_�F�*qA����6\�4�@�� �-jېI�q�������?B��#Ɵe�*|�÷�Wе !�`�(i3L�J)���� \L�1tSjv�����l��P��n�#�$a��o���H�RtV�^?�k�V�?����fJ��I����~uK7͍��|��W&":�ݚ�Н���w�w:�!�`�(i3�2�9�sye8�� scX{�X!,;�jmT�#Z�y��	�����u��r��!�`�(i3*�˜	����r"nCo��I�Ūe�ǩ"�4s2��ԜF��v��?���(1tSjv�!�`�(i3�Կ���p5��6V�|J���QE���(�o}��p>�!�!�`�(i3���%>�rGO�D mWN!�`�(i3��Ě�����}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ�c^����24���7�T�O�.�g3Z�)V��B�1'���5���s�s��M+�t�+!�`�(i3�g����&�P]�^qB���یHKz�Q��q��3���5�O�%E#P{y����M�V<�'������o�5�~NiQ3S����A��R�ߋ��V[ý��IX0F�MV�ҁGG�.Mm-;�C>��Ӛ��S�J\7Z$��k�4��x�S~p�A�W/��Wu�|#HK��A(�c���_G��Hb�8�u?��I!�`�(i3}�gv�oE�[��s�A>�xw'��M�v�����FK��|�H��4"�Կ���p5��6V�|��nF���<�W�.�P��=�ԇs�̢k���F�KD�Vr[/}>5��0�7<(�lb��� л��E�BS�+��U�,�P!6���r�����$XR�QܛOcOZail������&G!�`�(i3�����y��'����u��r��!�`�(i3�����n��)��RU��my$�N��o�/���;!�`�(i3.��fReU!�`�(i3����.��Ν�ʉ_��ݚ�Н��H�����������'����ݷ;���U;S����xQ�1tSjv�!�`�(i3�\>�ʘkN;LF�K�j�!�`�(i3�߆�p�h���/a�O����xQ�����@�ܵ�ҕ1�PS�B� �b��!�`�(i3�H��������P`��cG���`ö8�b(���sjߢiVr�r%)cA�C�)3vX�!�`�(i3A���P��6� ;h$	�(0f/-��8�b(���sjߢiVr�r%)cA�C�)3vX�!�`�(i3A���P��6� ;h$	���tY�:8�b(���sjߢiVr�r%)cA�C�)3vX�!�`�(i3�������l̲�2�!�n;�J���	��u�ܨ���@+�c�1ǺvK}� h�ҩ�!�`�(i3Q3S�����p��8��Lt���h�T�ns��m��B�_֭7.~t=� �!�`�(i3���F��O��ݚ�Н��Ra])n#��%O7G����:r���' �����%�gx{^4��*m!�`�(i3?�k�V�?����fJؔ�(�;giث���fJؚ�G�x )!�`�(i31���~!�`�(i3�G'�a@��6� ;h$	�W�L�sQ��|`��'��>�4Nu{ᵿ�����X� 2!�`�(i3��m�~r�DM3-���~�}��03p��|`��'��>�4Nu{ᵿ�����X� 2!�`�(i3��m�~r�D�Ÿ���H�}��03p��|`��'��>�4Nu{ᵿ�����X� 2!�`�(i3��O����k�r"nCo�A((���ڥ����A�}p���I
;Ȼs���ݚ�Н�!�`�(i3�Lt���h/��$�aZJ;_Q���Q�{;�X������I>������!�`�(i3���F��O��ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹���3�~\�0^˥�2��Z���/(_��)iƃ�;��|B���"�'�%d"�iF�a��ˀ�!e�ez8�US���W}V�U��)���Y;e�iKI/B޾Pb�i0[���S�J\7���_J��`L��Y-1ף�V�OnͶ�2��ibs��2[�a��o���zM#��m�!�`�(i3��4h�=Iz~r��V�n��dK�����fF0��hs�����F;p�	+��Q��:~Y&:��8�AԢ�a\�b7����"�A�;�֋`N��7�j2��9�,�n#,\ͨ܉p�u-/���y�8��C"��|U�O�-F}���V6w��EO"�̞��>���I�Ūe��Z�Y� (�6k�4d��Tٷ���
z�.�M�I����~u���P�|T����{7�R��ӟ-��ْ �%z�A�;�֋`N��7�j2��'Kb�|n���7���ө�O6�]Η^ś���k�i���ؠ��6���9�
z�.�MJ�A7��x��7���Zh|���!�`�(i3�I����~u���%��Y��k��^�1��dc�@c�����h�'�ɳ��<�6�Q=��ž�Ć�T���7X���c�}�:
��x�{�\��N�Ś�-����;�jmT�#Q���V�_�mS8<�n�ݚ�Н�|�au�(Z�H<�2�8��C"��E�g�������(ӈ���m�r����q�9�ͭ�M���V��+��Q��:~��/���bx���P�|T�T�����U(���B���ި���pj2�q�*t��}Dq�f����Mڷ�2v.^࣡N!�`�(i3iŞ�W�%3AԢ�a\�ɓ�~Ҡ	6d�dG�7:�R���Z�F�\Ȳ�r�r%)cA�%�\B�����x.�KnqQ������ݚ�Н��SSB������l�@�������įէ3��}Dq�f�N
������U�� ��!�`�(i3� ��U�_:��}Dq�f�8Uf[���!�`�(i3�L����j��W/�mƍ2���l�<�6�Q=��j�3����^�|ǔ����l���t�1C�G��HbH���!�`�(i3'-Bd8il�e���;X�W>�V��I�Ūe߰�	���1tSjv�!�`�(i3f���8�6�e���;���
`_�{_8�Y��=�}�Vݨ��}Dq�f�՝� s�#���k$ !�`�(i3��@h G0�H_��#��M��<̻�J�M���V��+��Q��:~�8w�B!�`�(i3���F��O�VA�ڦ�c4;�jmT�#��@h G0�H_��#��`����W��yM�5���%�+� h�ҩ�!�`�(i3졾�8 &F;p�	+��Q��:~�W�J��R��ӟ-���J��RQH�RtV�^!�`�(i3��=m緒Sr��3��ő��̼��nF���<�W�.�P�	��
�Q�}!�`�(i3�����!�`�(i3�B�'��a���p��b���ez8�US������`��kv޶Gl�e���;�z}+;��ݚ�Н�
�:qEp�;�P�t�5!�`�(i3$f��_Ub����pT�!�`�(i3'-Bd8il�e���;X�W>�V��I�Ūe߰�	���1tSjv�!�`�(i3QV�=��u:��_x�H_��#��O}�!��ƾ��7�j2��S]�_�_��u��r��!�`�(i3\���F�`y��Tٷ��N�$��+���a\Y�����J��RQH�RtV�^!�`�(i3���Mڷ�2v.^࣡N�I����~uK7͍��|��W&":�ݚ�Н�!�`�(i3�SSB������l�@�J��lb��j)����r^!�`�(i3�Ra])n#���r����!�`�(i3���Mڷ�2v.^࣡N�I����~u�5?�&P-�^��~_װs!�`�(i3!�`�(i3����E�El~pDa���̞J�2__���LefV�$����ݚ�Н�!�`�(i3���F��O�VA�ڦ�c4!�`�(i31���~!�`�(i3١w��zj�XYS��1��-P��C���c��b(�ԇ"'��&އ�L�Ģ�^r�r%)cA��gx�܈!�`�(i3HN��R��bP�63Z�t!�`�(i31���~!�`�(i3[�t��#�Β �r��1��-P�͹9^l4zױ��ԜF��iR$�Si"!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	����
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�\E�W��4b�^�#�n�i���w�6s���B�˭s;����_�� -]��V[ý��IX0F�MV�ҁGG�.Mm-;�d�G}%����3fGg��q�6��@�;��ʡ.>��'ž1�|�'����z.��W��!�`�(i3����j��3���B[=����e���A��s�R�b>3��g`
 ֢���@�k��}/ ���we��0�U+�qbp@�`
 ֢��.��� j�H]����j)����r^�]��W���Sd�[��q9+t�}b�0"qo�0�ʂ�j�Ï��	�l�lM�3 zM#��m����F�P�7��S��h��d\��H����o�γ�ha��o���H�RtV�^�I�K�B(�W ���t�1tSjv���6�����7*9uu!�`�(i3E�g�������(ӈ���m�r������6����Αk�]I	V��@��/�įէ3��}Dq�f�vx��c6���J��������;q��b+}y[՝� s�#���k$ �� л��Ԇo�	���q�ӘS��H����!�S_�_�mS8<�n�ݚ�Н�E�9�ؕ�^3rdS���I����~u���NM���!�`�(i3�2C9��o#�
z"H����t���m������� h�ҩ�!�`�(i3���D)��J�a$�Y dN�<@Iv��nt=:��:5A��p
�:qEp'{w#/ B!�`�(i3�G%�MP3�_~�:N��gKh���1�B.>!�`�(i3HN��R��bP�63Z�t!�`�(i35��
�4V��E9�}u��r��!�`�(i3i�]ʺ�
ǋ;�-mO�J�A7���ݚ�Н��Ra])n#5��
�4���ڌ�&-���x�'@�(��P�G�p�PXI����|�ݚ�Н���6����Αk�]I���,��~�B-�QŤ!�`�(i3�k��^�1̲�2�!��)��
�f��yM�B(p`D҉̖�7�j2����|��H�RtV�^!�`�(i3;+�'ն�%H=1b�ᅁ�:��!�`�(i3�̢k������D)����5������7���ө�)�F��3A�)Oq����ڽ�u� h�ҩ�!�`�(i3��|>�ğo���X��l8R��!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��jϤ�LǀP)���L��`����#Q���;�Ӏ�I:N�7�����t�T��?E-h��$^(?��"]�B���[:Fa�7��׏����Ļl�G�E�O�����"sS<�0�zG����ZAL�:!�`�(i3���y��lD�	Sz��
�GBQQY����#H�Yg�yi��v��BPlLO+��JתMܥ!�`�(i3'�^���������௴PJU���-|6�Ƃ)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0�7<(�lb����y��lD�7m�T��Ʈ+ˀa��z��2�,�$XR�QܛOcOZail������&G����l��P��n�#�$a��o���H�RtV�^�l\�6�'����7Z��n��뾦�!�`�(i3�e�MW���}�OCCfﾸb+}y[՝� s�#�=����T;�jmT�#�B�fL�ŋ;�-mO��ȭzB��6���9���H��R<z'�$쾹KK���������E�El~pDa��xR��\a%�G�&C�ez8�US�B�!����r�7���ө��i��o0��sOS���Z��oGM�о٫�Y�2]%�IG�p�P�➁q��^3ZiYX�m��Ӈk��fg�p5��Q��"��h��;��B� �b��!�`�(i3��s8��J�a$�Y ״$(�>g�!�`�(i3��jVѭ@!�`�(i3]a%ڔ�����;q��b+}y[!�`�(i3�5ߧE4��!�`�(i3�.2���	W��e5Z	�R/*__���Le<����t1tSjv�!�`�(i3*��^�"~HR�3]� *Ɋ��NM���
�:qEp'{w#/ B!�`�(i3�#�l+�����pƍ2���lĉ��%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j�_�Ƭ7~6O���N�ޓ;dE�\97*�SC&k@C�Ɨ0z�cUL��#R���2��2it��w�K�})9ͬ果��S�<Ԣ�7Z�:1�\mdЧ^{�j��$�'	���:<��j~�Q��g�]��`4Ƹ�$D@P�����g�I&�$a鯖U!dj`���=� ò'�����7y�	7�(�� ��S]ȋ�I���c�90��y�"v�W�Ep�_�d����\����z�5Y�IX0F�MV�ҁGG�.Mm-;�d�G}%����3f���K��M� ��l�J}�xjzӝ���I(͂�'�ɳ��!�`�(i3<�6�Q=��S<����K��!L��3w #�T�Z��&�2�����I��m�]�e���b���nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")z.��W����Q�Y�;y��v��\���
^�|#HK������ �'����u��r����#�a�Ą1 �u�.������&G!�`�(i3�)���IrŐ����l�K7͍��|��W&":�ݚ�Н���jVѭ@!�`�(i3�$|�ݲ�w&͏���M?��y�!�`�(i3q�\E��0d��ZS��o�]�S�*1�ó%2(!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�M��<:� �`�8j��M��%2�/�C���t�T��?E-h��$^(?��"]�B���[:Fa�7�����~�Ln�cqgF}�P�|�bs��2[�a��o���zM#��m�!�`�(i3��4h�=Iz~r��V�n��dK�����fF0��hs�����n��0�5	x!�`�(i3/ ���we��0�U+�qbp@��'��o�u:��_x25���w����;q�{_8�Y��=�}�Vݨ��}Dq�f�/N2~-��x�f7﹏!�`�(i3%��v�ڹ߆�p�h��d��JXl'�T��~��?u��C@!�`�(i3.�
9� ���(ٗ.;���JTv�䵶
�t��T&��ۥ`�M?��y�!�`�(i3�!AaiT��G��Hb� h�ҩλ�(1l�jG���Z��o!�`�(i3E�g�������(ӈ���m�r����B�'��a���p��b��L,d\P��n��>�my$�N��o�/���;!�`�(i3�w[��r^�/;�������I����~u/��kOT�Ra])n#���r����hs�����n��0�5	x!�`�(i3s���IK^�!��w��1�ó%2(!�`�(i3�$|�ݲ��'����u��r��!�`�(i3�kv޶Gl���m\g�Y��0:�rs�i�E�8�w��ӭu:��_x�H_��#���QtόH�i!�`�(i3�5ߧE4��!�`�(i3e��4&�N��r�������;qu�#:I�˜!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�MТKH�{?ۄQ�0g��L�Y}śT嫞ic)�̩�'��N��v�8�u?��I� ��U�_:_f.�}�ٷx�Z��x�́���y�I��Mq��+����$��m�4VG���D)��+c��p*OZ鎬�������(������P`����^�"�B��\��[��&k@C�Ɨ0z�cUL0:_\�c�XYS����u'��W-37�˱�5ఽ��`g�]C�����i#���ϸ��#|S������3[�u8��v1a{J�^�|n�M�!�`�(i3!�`�(i3J�]�RU�`�����hy�/B/���^!�������>)�ak�m6!�`�(i3,54��]��)�4!�,�ttT�r�pΚ�w]��Ɋ]�!�`�(i3�&8�,������k�v2<�����h�? "a��Q�V!�(�!�`�(i3�X;p`�V�׍A�f�?ǉ�=��<E�f��V�mK�b6�X�$�!�`�(i3�;�����^��&X!=�t����}�(�
4��c��^�
E��#	����J!�`�(i3r�(���i�lK�f�?ǉ�=?�ᒹ�G�!�`�(i3!�`�(i3!�`�(i3��\��,&߰��U��f�?ǉ�=���gRI/)�ak�m6!�`�(i3!�`�(i3���Z�N�j����t���hQ�GvE�<�W������!�`�(i3!�`�(i3-���i�4(��i缔]���W����L�z��̾_4k&}ǝ^3!�`�(i3!�`�(i3HƏ~g��ղT�D3H	hDJ��3Y� 2��4����7
!�`�(i3!�`�(i36�ŏ ���N���B
���������b�Xϋ?@,�Xʚ@h!�`�(i3!�`�(i3fC��T����ܼ�_`Ogkl@`��m'��r�Nt[NzigzA=v)-��,ufOX�mCf�?ǉ�={p�R�I8$vVqYY!�`�(i3!�`�(i3J�]�RU�`����y��j��k��V��e�LtW��e���d�tAAI�O����0 �;t��I���yR���/�"����0@�pgd@!�`�(i3!�`�(i3!�`�(i3��P��fn�[q�<i缔]���7p�J��PW�o#�_T��!�`�(i3!�`�(i3!�`�(i38~<�o�?��bTg�zϾZ��s?�t}~�Y���(���;����f!�`�(i3!�`�(i3!�`�(i3�F�7��Y�
�cc�V�/�"����0�:C&e�!�`�(i3!�`�(i3!�`�(i3���u�UgF˯�+)��&�C�/�#�@�o0�&�v�x!�`�(i3!�`�(i3/;�Ly�A<���O�0��s���4@Q�/���hy�_�⥳�"_!�`�(i3!�`�(i3!�`�(i3�9�x��/�"���꤭%�3��{!�`�(i3!�`�(i3!�`�(i3�X�w���A�:JϮ�M?�_�9�!�`�(i3!�`�(i3!�`�(i3�X;p`�l.�	�C�Y��j3���k��0H!�`�(i3!�`�(i3!�`�(i3���*[UxGZt%��m&<g+b󆤐=!�`�(i3!�`�(i3!�`�(i3С���?�1 `m|V��������iA'R�	!�`�(i3!�`�(i3!�`�(i3�n�a#��E��\��[��f�?ǉ�=���L��T!�`�(i3!�`�(i3!�`�(i3@�m��nmv�:����TBd��p!�`�(i3!�`�(i3!�`�(i3�X;p`���C�,�4G�E
b�+|!�`�(i3!�`�(i3!�`�(i3!�`�(i3��n�T���v��X�<�!�d�<p�m����v{��lw	�Kk
�&1<5F��e�R�CB���+����$�o��A�3~9�W6�b�˱�h�Vy�