��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S��������ߪD?=N��J��S������!P7TǱ�J���G�J6�qQ��iQ�����-v�ZN��pV�!���}��J6�qQ��J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag����pH��q$.:&R�nU���T��ײ2��>���^k�/7�?1�(�c��ߘ�]��|�G��f�:��#tC��o�Rb�v �mD�?�D��L���_�L�Ȳ�V�溜��D�,�H�9� I�����5O|��N�w	*D���y&�f��+K��[y��ڂFWe5)�o_ ������/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�7Y[���G���d�֗r�5�c$e
�9��Ax!P����yџY{P�h$�;��I���*�F�l����Iݱ�.���� �bRw�����IL�+�{Dr[���Ѹ�t����g�*�$}����L�v&�2��߶�5��1y�HU��GAݐ_�!����P�>��H3NVI۷� �{K��"\����v�����V+�9ުE,?����>�8p��Z~G0�M6w���8Ǎѻ�%�R(�h�J�yU�k�.
���dt�{������K�䒆	�_3�3k����tċ^9t��M�����=T��i��B�����$b�[��|�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯�^��N�&��?�2�1p�r���q P�^�&d�A|?_W�\I��^�َ2V�N�u�k1i�f1?�نN��_�Q�L���E����[�/�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_E$ô&y��aC�h�>�N{a�9Ow�Y��k��ı��*���q{?d']la�b����M:��;6aJVlO/2>� zM흜5���_M	������Q�^�y�zL͊�q�����$�!h��6h�烋l�;�w����g�&�0m�b9���:&�>��s�䉌�+B4��ղ�^yP��b�G�lnO���t�S+ɭ(��
��,ysA�U�y�S�ŇO�[l���8l@U}�8���[��C��!�`�(i3�E����F���8�TP����������s	IB�;�5�}�]���!�`�(i3зq8�Ј)w�<�_N$��)bX����<7e �Ç�t�<H�W�h���Q�#<4^�!�`�(i3v�ј�"��Z鎬���������o�	Ql��ɐ!�`�(i3N�By3��<�]�!��5��E0�b��8�#e۽V��*J !�`�(i3N�By3��<�]�!����M[��Ǣ�˩��*��!�`�(i3�����5	���]���>����C��x��� ��2�w���������e.��xu	���S8�bM� 2)G��8���/��P���w�m���d�!�`�(i3v�ј�"��Z鎬�����	�7 �#�iK�D�b=| ���jN�By3��<�]�!����M[��Ǣ+���G��!�`�(i3�����5	���]���>����CΤ��8�%Y�����U�����E��@IE�U��>��l%i�-I����hoDy����g-C�#��R7G#+��\w��0](@X~�H:���������03R���TD���rs�i���	�>�g��U-�e�,���6+�����0��G��e���������t�SI��w��,>����CΊE\r���!�`�(i3�����E��@IE�U��>��l%i�-���s�`�zM#��m��E����F��j���0z�cULm�Y�ڱ��5���_M	"j���b7|#9���EOJ�uxm�Ww3i�|�"�,�>E���TD���rs�i��;m��"xd#���>��CyW�f�tR�wX���Y�_�����!��R-!�`�(i3��(�
t�������2%=dϖ�i�!�B����� j���tN2s��/~.)��3\�R�F*}�c}��uO�b�^��\/ɭ��:�Q��ņD^�NË�����8�9Ѽã� Oag��Ц��#�"�Q:�{�1k�ZV"���:��#tC���,?a��Q\�_qť��[�޿3ų�̿}�
�?�	�%��6�1�#��d_зq8�Ј'���Xw�%G��lyl������!�`�(i3!�`�(i37s�9���o>��l%i�-5�e`��9S�n�(�a_1�f�����Q]� _ό���.�}�
�?���)�δ��+�qy�t4��_���'���Xw���,D�H�p0�����dܟz�3l;X��]�!����w�Հ�b02�ORR6��-z!�`�(i37s�9���o>��l%i�-�u��Y'Gish�Ž�Լ^=Г�m��Jn,���`ό���.�}�
�?��W�3�-[)��V���зq8�Ј'���Xw���,D|�|��f3�Y$�J��;"�,�>E���]�!��ߞ��-���L5ӥ���������p�PB����A�����]o{�k?���ʟ�DFV�t%>^����80�i�!�`�(i3Y%T��BP	�I]����.�Ӂv�u�o�\�A�|P;៪p�:����I8I����T@a��F�!�O��1���Sns&����rS�h���^.�]�YǯXan��o��pL5ӥ���b�W1c�͌�Nf����t%>^��?�y��hL5ӥ����B��+ H7�ܥ��2��T��o�B�t%>^��?�y��hL5ӥ���d��P���lC��ۺ_~�x��+�`:�H/��$���� ��\��+0�NҰ�y)���y���7m�!t?' t����/�nrm؊(��dט�w��׺8|MW���0o�_o�7�ܥ��2��P:q�hg�4�+/r��bQK����0�VC �7)N�J�wII��'��vbëdP���|�r�HzL͊�q�����cj%������4��k�y'��a[��gAQ+��t��h~�,��E���Q]� _ό���.�}�
�?�#l'U:�g[-�¾L���d�٣���N N�S��E �����VF�˷�]+W��L��'���Xw���,DFmғO�4}~n���,a�n`5�fK�\w��0]b!��uፊ5�j�))O�LYw9���]�!����w�Հ��a�e56<, �c��β��+�J���q���U��@����gG|�w��DKCϗ(���7s�9���o>��l%i�-He�-�c��d��]�Q�}J�AZ鎬�������(����F�dHP����|�J!b%�ZV���"X��[��Q[R�7He�-�c��3E M0�F�T��BZ鎬����Y�V��#q���`����C�%�_�S�
ut�q���U�`V�-(�e<�ߢěf%װ$��_�zM#��m�{�R�$�V�<�xwu�P�#c8o7C?���f��3ALaX��T.�D%��Ai_�ܛ%w�*�7�����'[�q{��xR�rf����˻*���J=��N6�;�c�uU�,r�-!�`�(i3�%5�����Wo���˃�e�����Wo���˃lp�h1���	;	�J����q�U�%t̓�@�H�\�{\��xA�[���D����/y��$ŧ��3o��~��U�WF8юn:�Q��?�\���>�(��G rgA�iK�D�b=��p�:�F!��D�����k$ !�`�(i3!�`�(i3Р�(�V���e�Ѧ֯���,--�O��Ud�^F�)�u]�MP��(R\֎u�D��u�(nP?��!��4���~�I��-��R>ݒ��liF��ê�\���S)��p�:�F!��D�����k$ !�`�(i3!�`�(i3٪�o�_&��E\r�������;q��)�δ��1�ak-�v�?�{�,�+����$�� 0�Z����Wj4�O	����C�(R\֎u�D��u�(n�s*�4��A��U�[�m��U��)���Y;e�iK-pm!9�>ֱ�q��,��ur�5p�T�ۣ�� L�>�0z�cULA6{'8�0��9gP�U,��!:����Г8���/�D,�n�G���rN�>�YS
?s�����W�0I��uy�_$��V�{y����i�q,?5qr4�Ў���<�e��BF�U���e��d9=���u��r��;[�T����	;	�J��f�Ϡ�����b+}y[�D�����O����&{�Iћ<��%��v���#�-�p��5p�T�ۺ��7Z��q(����b�z'hۉ)��d�7�qā��̰�!�Xy|�W�(�[�*%��v���#�-�p���p�:�!�`�(i3��$�\%e��}Dq�f�o;�Ul�|�Ƀ�?PAn�#�7�;�j)����r^*qA����6\�4�@�� �-j�1tSjv��V�qZ%	R>ݒ��lĪN�!Z�������	;	�J�����I-�X�7���������U���g��%5�������p1��#�-�p��5p�T�ۺ��7Z��w{���@�ّJ8��e��2
-�����9gUS����a$�/=7�7K�PO`�� \)�(R\֎u�D��u�(na��[%���K�&�a��+���q���i+��_1�f���!�`�(i3]
���7ϥ���WՁ��̰�!i�q8�2t�ݡ��1������$~@�J�g�*~,�H�͛���Ě�����ˣ�X7,R��(�ٰ�Ř�hsGS��c��ّJ8��e��2
-���������=��߸��S�Ȍp�M���)~A�\MU��$ϙRl�b�Qx�v�^�����8^�Xe�)զޢ:ͤ�B@����=�?@o�7qz+�XЙMǿI?��^�r-XgJ,�|d�n���G΂�M�{�|L�.r�$����#o�]�ʄ�v�4�?zmU�WF8юn�jjC�_�vާ���虾�b+}y[���$A ���U�E�u�N�iK�D�b=��p�:�F!��D��M����ge�����'�ekl������a�h&�,\ަ�It��+g[�DsQ�V�r[��7�y&��˼S����#X荂:\�C4%̈́�A��4�h���6X�Obq0�~����O�΃S�������௴PJU��ĤI�v�����&8�,�e'M�)�p�_��SW86�όz#�<ո1_�
774\51�]2�t��MJT��
!�7�R�"�*}�r������&Ve�!�`�(i3�X;p`�!͙��04n$v��a����^=�0y��bm�ms�����I�[�ȫw��`U@!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�0�����nX:��+�k_����Zv���;-����`�����uk�3��H9�r����ؾ<k�[��x�ܽ���X;p`�T���'/�>�r����`�4,�pI�!�`�(i3�X;p`���.�ֽ�f�?ǉ�=��5@~Ju*k`Ë��!�`�(i3��*�{6�
�cc�V�S7�8�8}�� �с�'(�U�c�&8�,��
�Q!}-[��u�����NPB7Ԅ���V��(��sW��|E�q��w\F�k S���zǣ©���>�@�C5]�꼧5#b|���Mk S���zǣ©�� ��ߕ!�`�(i3!�`�(i3�G8T�w�n;���C#����d�E����'m�|g�~p!ۓ<���O�0��s���4@Q�/�r�VU���l����S�U젩`#36��T�%G�͚���v�h̤�Vl����STl�����)��.��f�?ǉ�=եa������X;p`�(�����Y�ay}M�!�`�(i3U�%
�b9�?|�i�Y�#�m⇗&8�,�j%a}�C})�^�\
���&~^)�&8�,�cop ���6�G|��� ���)�{� �"czZ�����
�%���F{/�����,([�y����ŕ-�Щ��O�*���]�ܯ���@Tvs�!�`�(i3�$�~c/�R��ŭ�.���ߠ����9
4�٩S��I�����Y>�څI������M�Mb�:u�!����3���3E M0�~�O������ԕaOf���x�f7﹏S��I���f�E�7��J~��u�'��۬�vDvA#&��Q-�b�+�